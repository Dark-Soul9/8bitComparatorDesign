magic
tech sky130A
magscale 1 2
timestamp 1685814321
<< checkpaint >>
rect -3932 -3932 16985 19129
<< viali >>
rect 1501 12393 1535 12427
rect 4077 12393 4111 12427
rect 5365 12393 5399 12427
rect 8493 12393 8527 12427
rect 10241 12393 10275 12427
rect 2513 12325 2547 12359
rect 7757 12325 7791 12359
rect 8401 12325 8435 12359
rect 2053 12189 2087 12223
rect 2329 12189 2363 12223
rect 2697 12189 2731 12223
rect 4353 12189 4387 12223
rect 6561 12189 6595 12223
rect 7481 12189 7515 12223
rect 8125 12189 8159 12223
rect 8677 12189 8711 12223
rect 9137 12189 9171 12223
rect 10609 12189 10643 12223
rect 1777 12121 1811 12155
rect 2237 12121 2271 12155
rect 5641 12121 5675 12155
rect 8401 12121 8435 12155
rect 9965 12121 9999 12155
rect 2881 12053 2915 12087
rect 6745 12053 6779 12087
rect 7941 12053 7975 12087
rect 8217 12053 8251 12087
rect 9321 12053 9355 12087
rect 10517 12053 10551 12087
rect 10333 11849 10367 11883
rect 5549 11781 5583 11815
rect 11345 11781 11379 11815
rect 1409 11713 1443 11747
rect 3525 11713 3559 11747
rect 4077 11713 4111 11747
rect 4629 11713 4663 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 7941 11713 7975 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 9137 11713 9171 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 10977 11713 11011 11747
rect 1777 11645 1811 11679
rect 3617 11645 3651 11679
rect 4169 11645 4203 11679
rect 6009 11645 6043 11679
rect 7757 11645 7791 11679
rect 8677 11645 8711 11679
rect 2053 11577 2087 11611
rect 3065 11577 3099 11611
rect 5825 11577 5859 11611
rect 8033 11577 8067 11611
rect 10609 11577 10643 11611
rect 1593 11509 1627 11543
rect 2237 11509 2271 11543
rect 3341 11509 3375 11543
rect 3985 11509 4019 11543
rect 4445 11509 4479 11543
rect 6377 11509 6411 11543
rect 7573 11509 7607 11543
rect 9045 11509 9079 11543
rect 1685 11305 1719 11339
rect 2329 11305 2363 11339
rect 4445 11305 4479 11339
rect 10333 11305 10367 11339
rect 10793 11305 10827 11339
rect 1961 11237 1995 11271
rect 2513 11237 2547 11271
rect 4997 11237 5031 11271
rect 5641 11237 5675 11271
rect 9965 11237 9999 11271
rect 11345 11237 11379 11271
rect 3433 11169 3467 11203
rect 3893 11169 3927 11203
rect 5733 11169 5767 11203
rect 10977 11169 11011 11203
rect 1409 11101 1443 11135
rect 2789 11101 2823 11135
rect 3065 11101 3099 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 5181 11101 5215 11135
rect 5273 11101 5307 11135
rect 7113 11101 7147 11135
rect 7481 11101 7515 11135
rect 7665 11101 7699 11135
rect 8033 11101 8067 11135
rect 8769 11101 8803 11135
rect 9689 11101 9723 11135
rect 9781 11101 9815 11135
rect 10057 11101 10091 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10885 11101 10919 11135
rect 11069 11101 11103 11135
rect 11529 11101 11563 11135
rect 3801 11033 3835 11067
rect 4261 11033 4295 11067
rect 4813 11033 4847 11067
rect 4997 11033 5031 11067
rect 6101 11033 6135 11067
rect 6837 11033 6871 11067
rect 9505 11033 9539 11067
rect 10793 11033 10827 11067
rect 1869 10965 1903 10999
rect 2329 10965 2363 10999
rect 2881 10965 2915 10999
rect 3249 10965 3283 10999
rect 2053 10761 2087 10795
rect 2421 10761 2455 10795
rect 2973 10761 3007 10795
rect 7941 10761 7975 10795
rect 10149 10761 10183 10795
rect 2789 10693 2823 10727
rect 5825 10693 5859 10727
rect 7297 10693 7331 10727
rect 8277 10693 8311 10727
rect 8493 10693 8527 10727
rect 9689 10693 9723 10727
rect 11253 10693 11287 10727
rect 1409 10625 1443 10659
rect 1961 10625 1995 10659
rect 2237 10625 2271 10659
rect 6193 10625 6227 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 7573 10625 7607 10659
rect 8033 10625 8067 10659
rect 6009 10557 6043 10591
rect 6377 10557 6411 10591
rect 7757 10557 7791 10591
rect 10241 10557 10275 10591
rect 10701 10557 10735 10591
rect 3157 10489 3191 10523
rect 6469 10489 6503 10523
rect 7665 10489 7699 10523
rect 10057 10489 10091 10523
rect 10517 10489 10551 10523
rect 10793 10489 10827 10523
rect 10885 10489 10919 10523
rect 1593 10421 1627 10455
rect 2973 10421 3007 10455
rect 6009 10421 6043 10455
rect 6101 10421 6135 10455
rect 6929 10421 6963 10455
rect 8125 10421 8159 10455
rect 8309 10421 8343 10455
rect 4721 10217 4755 10251
rect 5641 10217 5675 10251
rect 7665 10217 7699 10251
rect 10517 10217 10551 10251
rect 10333 10149 10367 10183
rect 11345 10149 11379 10183
rect 1961 10081 1995 10115
rect 1409 10013 1443 10047
rect 1869 10013 1903 10047
rect 2145 10013 2179 10047
rect 2789 10013 2823 10047
rect 3157 10013 3191 10047
rect 3341 10013 3375 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 4537 10013 4571 10047
rect 5089 10013 5123 10047
rect 5457 10013 5491 10047
rect 7389 10013 7423 10047
rect 8217 10013 8251 10047
rect 11529 10013 11563 10047
rect 3525 9945 3559 9979
rect 4445 9945 4479 9979
rect 5273 9945 5307 9979
rect 5365 9945 5399 9979
rect 7481 9945 7515 9979
rect 7697 9945 7731 9979
rect 10057 9945 10091 9979
rect 1593 9877 1627 9911
rect 7205 9877 7239 9911
rect 7849 9877 7883 9911
rect 8033 9877 8067 9911
rect 4813 9605 4847 9639
rect 5917 9605 5951 9639
rect 1777 9537 1811 9571
rect 2329 9537 2363 9571
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 4261 9537 4295 9571
rect 4537 9537 4571 9571
rect 4629 9537 4663 9571
rect 5733 9537 5767 9571
rect 5825 9537 5859 9571
rect 6101 9537 6135 9571
rect 6193 9537 6227 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7573 9537 7607 9571
rect 7849 9537 7883 9571
rect 8309 9537 8343 9571
rect 8585 9537 8619 9571
rect 8953 9537 8987 9571
rect 9045 9537 9079 9571
rect 10149 9537 10183 9571
rect 6377 9469 6411 9503
rect 6745 9469 6779 9503
rect 7665 9469 7699 9503
rect 8125 9469 8159 9503
rect 3709 9401 3743 9435
rect 7757 9401 7791 9435
rect 8493 9401 8527 9435
rect 1869 9333 1903 9367
rect 2237 9333 2271 9367
rect 2421 9333 2455 9367
rect 3525 9333 3559 9367
rect 4353 9333 4387 9367
rect 5549 9333 5583 9367
rect 8033 9333 8067 9367
rect 8677 9333 8711 9367
rect 8953 9333 8987 9367
rect 10333 9333 10367 9367
rect 10609 9333 10643 9367
rect 5089 9129 5123 9163
rect 9045 9129 9079 9163
rect 2513 9061 2547 9095
rect 8217 9061 8251 9095
rect 10057 9061 10091 9095
rect 2237 8993 2271 9027
rect 2881 8993 2915 9027
rect 8309 8993 8343 9027
rect 9413 8993 9447 9027
rect 10241 8993 10275 9027
rect 2789 8925 2823 8959
rect 5457 8925 5491 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 8125 8925 8159 8959
rect 8401 8925 8435 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 10333 8925 10367 8959
rect 10481 8925 10515 8959
rect 10798 8925 10832 8959
rect 4905 8857 4939 8891
rect 9781 8857 9815 8891
rect 10609 8857 10643 8891
rect 10701 8857 10735 8891
rect 5105 8789 5139 8823
rect 5273 8789 5307 8823
rect 7941 8789 7975 8823
rect 10977 8789 11011 8823
rect 1593 8585 1627 8619
rect 9571 8585 9605 8619
rect 10333 8585 10367 8619
rect 11253 8585 11287 8619
rect 2329 8517 2363 8551
rect 2697 8517 2731 8551
rect 5549 8517 5583 8551
rect 9321 8517 9355 8551
rect 9781 8517 9815 8551
rect 11069 8517 11103 8551
rect 1409 8449 1443 8483
rect 2605 8449 2639 8483
rect 2789 8449 2823 8483
rect 3157 8449 3191 8483
rect 3341 8449 3375 8483
rect 3433 8449 3467 8483
rect 3709 8449 3743 8483
rect 4537 8449 4571 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 5365 8449 5399 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 6009 8449 6043 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7389 8449 7423 8483
rect 9045 8449 9079 8483
rect 9137 8449 9171 8483
rect 9873 8449 9907 8483
rect 10425 8449 10459 8483
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 3065 8381 3099 8415
rect 3525 8381 3559 8415
rect 4445 8381 4479 8415
rect 6193 8381 6227 8415
rect 7665 8381 7699 8415
rect 3893 8313 3927 8347
rect 5181 8313 5215 8347
rect 9413 8313 9447 8347
rect 11069 8313 11103 8347
rect 2973 8245 3007 8279
rect 5733 8245 5767 8279
rect 6929 8245 6963 8279
rect 7205 8245 7239 8279
rect 7573 8245 7607 8279
rect 9321 8245 9355 8279
rect 9597 8245 9631 8279
rect 9965 8245 9999 8279
rect 10517 8245 10551 8279
rect 1685 8041 1719 8075
rect 2697 8041 2731 8075
rect 4077 8041 4111 8075
rect 4261 8041 4295 8075
rect 6101 8041 6135 8075
rect 9597 8041 9631 8075
rect 3249 7973 3283 8007
rect 5273 7973 5307 8007
rect 6469 7973 6503 8007
rect 7481 7973 7515 8007
rect 8677 7973 8711 8007
rect 9229 7973 9263 8007
rect 9321 7973 9355 8007
rect 11345 7973 11379 8007
rect 6561 7905 6595 7939
rect 7113 7905 7147 7939
rect 7573 7905 7607 7939
rect 8769 7905 8803 7939
rect 9689 7905 9723 7939
rect 1961 7837 1995 7871
rect 2053 7837 2087 7871
rect 2201 7837 2235 7871
rect 2421 7837 2455 7871
rect 2559 7837 2593 7871
rect 2973 7837 3007 7871
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 3617 7837 3651 7871
rect 3893 7837 3927 7871
rect 3985 7837 4019 7871
rect 4537 7837 4571 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 6285 7837 6319 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 11529 7837 11563 7871
rect 2329 7769 2363 7803
rect 2789 7769 2823 7803
rect 5273 7769 5307 7803
rect 1501 7701 1535 7735
rect 3525 7701 3559 7735
rect 4445 7701 4479 7735
rect 8217 7701 8251 7735
rect 8953 7701 8987 7735
rect 9965 7701 9999 7735
rect 2237 7497 2271 7531
rect 2881 7497 2915 7531
rect 5381 7497 5415 7531
rect 7297 7497 7331 7531
rect 5181 7429 5215 7463
rect 7665 7429 7699 7463
rect 1409 7361 1443 7395
rect 2789 7361 2823 7395
rect 3065 7361 3099 7395
rect 3157 7361 3191 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 7481 7361 7515 7395
rect 7573 7361 7607 7395
rect 7849 7361 7883 7395
rect 11253 7361 11287 7395
rect 1777 7293 1811 7327
rect 2329 7293 2363 7327
rect 2145 7225 2179 7259
rect 1593 7157 1627 7191
rect 2697 7157 2731 7191
rect 3801 7157 3835 7191
rect 3985 7157 4019 7191
rect 5365 7157 5399 7191
rect 5549 7157 5583 7191
rect 10977 7157 11011 7191
rect 3893 6953 3927 6987
rect 4537 6953 4571 6987
rect 9229 6953 9263 6987
rect 11069 6953 11103 6987
rect 5181 6885 5215 6919
rect 5549 6885 5583 6919
rect 10241 6885 10275 6919
rect 3893 6817 3927 6851
rect 11253 6817 11287 6851
rect 3801 6749 3835 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 9045 6749 9079 6783
rect 9229 6749 9263 6783
rect 9965 6749 9999 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 4353 6681 4387 6715
rect 4558 6681 4592 6715
rect 10701 6681 10735 6715
rect 10793 6681 10827 6715
rect 4169 6613 4203 6647
rect 4721 6613 4755 6647
rect 4813 6613 4847 6647
rect 9413 6613 9447 6647
rect 10057 6613 10091 6647
rect 4537 6409 4571 6443
rect 8125 6409 8159 6443
rect 10977 6409 11011 6443
rect 7021 6341 7055 6375
rect 7237 6341 7271 6375
rect 7757 6341 7791 6375
rect 7849 6341 7883 6375
rect 8401 6341 8435 6375
rect 10425 6341 10459 6375
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 5273 6273 5307 6307
rect 5365 6273 5399 6307
rect 5825 6273 5859 6307
rect 5917 6273 5951 6307
rect 6101 6273 6135 6307
rect 7665 6273 7699 6307
rect 8304 6273 8338 6307
rect 8493 6273 8527 6307
rect 8676 6273 8710 6307
rect 8769 6273 8803 6307
rect 9505 6273 9539 6307
rect 9781 6273 9815 6307
rect 10333 6273 10367 6307
rect 10517 6273 10551 6307
rect 10701 6273 10735 6307
rect 10793 6273 10827 6307
rect 11069 6273 11103 6307
rect 2697 6205 2731 6239
rect 5641 6205 5675 6239
rect 5733 6205 5767 6239
rect 8033 6205 8067 6239
rect 6101 6137 6135 6171
rect 7481 6137 7515 6171
rect 9597 6137 9631 6171
rect 9689 6137 9723 6171
rect 10793 6137 10827 6171
rect 5089 6069 5123 6103
rect 7205 6069 7239 6103
rect 7389 6069 7423 6103
rect 9321 6069 9355 6103
rect 10149 6069 10183 6103
rect 6193 5865 6227 5899
rect 9781 5865 9815 5899
rect 9965 5865 9999 5899
rect 10885 5865 10919 5899
rect 5641 5797 5675 5831
rect 11345 5797 11379 5831
rect 1409 5729 1443 5763
rect 3433 5729 3467 5763
rect 6469 5729 6503 5763
rect 7941 5729 7975 5763
rect 5457 5661 5491 5695
rect 5549 5661 5583 5695
rect 5733 5661 5767 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 6653 5661 6687 5695
rect 7113 5661 7147 5695
rect 7205 5661 7239 5695
rect 7481 5661 7515 5695
rect 7665 5661 7699 5695
rect 8033 5661 8067 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 11529 5661 11563 5695
rect 3157 5593 3191 5627
rect 6837 5593 6871 5627
rect 9933 5593 9967 5627
rect 10149 5593 10183 5627
rect 5917 5525 5951 5559
rect 7021 5525 7055 5559
rect 7389 5525 7423 5559
rect 10609 5525 10643 5559
rect 7849 5321 7883 5355
rect 1409 5253 1443 5287
rect 1777 5253 1811 5287
rect 4445 5253 4479 5287
rect 5733 5253 5767 5287
rect 5825 5253 5859 5287
rect 7481 5253 7515 5287
rect 7573 5253 7607 5287
rect 8217 5253 8251 5287
rect 2421 5185 2455 5219
rect 5636 5185 5670 5219
rect 6008 5185 6042 5219
rect 6101 5185 6135 5219
rect 7389 5185 7423 5219
rect 7987 5185 8021 5219
rect 8125 5185 8159 5219
rect 8400 5185 8434 5219
rect 8493 5185 8527 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 10425 5185 10459 5219
rect 11345 5185 11379 5219
rect 2697 5117 2731 5151
rect 8677 5117 8711 5151
rect 7205 5049 7239 5083
rect 7757 5049 7791 5083
rect 5457 4981 5491 5015
rect 10517 4981 10551 5015
rect 11161 4981 11195 5015
rect 1856 4777 1890 4811
rect 5089 4777 5123 4811
rect 10057 4777 10091 4811
rect 1593 4641 1627 4675
rect 10977 4641 11011 4675
rect 5641 4573 5675 4607
rect 5779 4573 5813 4607
rect 5871 4573 5905 4607
rect 6145 4573 6179 4607
rect 7665 4573 7699 4607
rect 7813 4573 7847 4607
rect 8171 4573 8205 4607
rect 10149 4573 10183 4607
rect 10425 4573 10459 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 11253 4573 11287 4607
rect 3617 4505 3651 4539
rect 3801 4505 3835 4539
rect 6006 4505 6040 4539
rect 7941 4505 7975 4539
rect 8033 4505 8067 4539
rect 10517 4505 10551 4539
rect 10609 4505 10643 4539
rect 6285 4437 6319 4471
rect 8309 4437 8343 4471
rect 10241 4437 10275 4471
rect 11437 4437 11471 4471
rect 5733 4233 5767 4267
rect 7665 4233 7699 4267
rect 8033 4165 8067 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 2421 4097 2455 4131
rect 4445 4097 4479 4131
rect 4537 4097 4571 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 5549 4097 5583 4131
rect 5825 4097 5859 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 7805 4097 7839 4131
rect 7941 4097 7975 4131
rect 8161 4097 8195 4131
rect 8309 4097 8343 4131
rect 9413 4097 9447 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 10517 4097 10551 4131
rect 11253 4097 11287 4131
rect 2697 4029 2731 4063
rect 5181 4029 5215 4063
rect 9873 4029 9907 4063
rect 10241 4029 10275 4063
rect 10333 4029 10367 4063
rect 10793 4029 10827 4063
rect 1593 3961 1627 3995
rect 1869 3961 1903 3995
rect 10977 3961 11011 3995
rect 4721 3893 4755 3927
rect 9689 3893 9723 3927
rect 10701 3893 10735 3927
rect 5567 3689 5601 3723
rect 8677 3689 8711 3723
rect 9137 3689 9171 3723
rect 10241 3689 10275 3723
rect 9413 3621 9447 3655
rect 1593 3553 1627 3587
rect 3341 3553 3375 3587
rect 3617 3553 3651 3587
rect 5825 3553 5859 3587
rect 6561 3553 6595 3587
rect 7849 3553 7883 3587
rect 8217 3553 8251 3587
rect 8493 3553 8527 3587
rect 9045 3553 9079 3587
rect 10425 3553 10459 3587
rect 3801 3485 3835 3519
rect 5917 3485 5951 3519
rect 6377 3485 6411 3519
rect 6469 3485 6503 3519
rect 6745 3485 6779 3519
rect 6835 3485 6869 3519
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 7481 3485 7515 3519
rect 7941 3485 7975 3519
rect 8769 3485 8803 3519
rect 9229 3485 9263 3519
rect 10149 3485 10183 3519
rect 6285 3417 6319 3451
rect 7389 3417 7423 3451
rect 8953 3417 8987 3451
rect 6009 3349 6043 3383
rect 7021 3349 7055 3383
rect 7665 3349 7699 3383
rect 10425 3349 10459 3383
rect 1777 3145 1811 3179
rect 4629 3145 4663 3179
rect 4905 3145 4939 3179
rect 5457 3145 5491 3179
rect 6009 3145 6043 3179
rect 8861 3145 8895 3179
rect 9965 3145 9999 3179
rect 10885 3145 10919 3179
rect 11161 3145 11195 3179
rect 2421 3077 2455 3111
rect 5181 3077 5215 3111
rect 6929 3077 6963 3111
rect 7941 3077 7975 3111
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5273 3009 5307 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 5641 3009 5675 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 6745 3009 6779 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 7713 3009 7747 3043
rect 7849 3009 7883 3043
rect 8124 3009 8158 3043
rect 8217 3009 8251 3043
rect 8768 3009 8802 3043
rect 9505 3009 9539 3043
rect 10793 3009 10827 3043
rect 11345 3009 11379 3043
rect 4169 2941 4203 2975
rect 4445 2941 4479 2975
rect 5733 2941 5767 2975
rect 8309 2941 8343 2975
rect 8401 2941 8435 2975
rect 2329 2873 2363 2907
rect 6469 2873 6503 2907
rect 9781 2873 9815 2907
rect 2053 2805 2087 2839
rect 7205 2805 7239 2839
rect 7573 2805 7607 2839
rect 6009 2601 6043 2635
rect 7849 2601 7883 2635
rect 10425 2601 10459 2635
rect 10885 2601 10919 2635
rect 11161 2601 11195 2635
rect 5825 2533 5859 2567
rect 10149 2533 10183 2567
rect 1409 2465 1443 2499
rect 3433 2465 3467 2499
rect 5457 2465 5491 2499
rect 7481 2465 7515 2499
rect 3801 2397 3835 2431
rect 5641 2397 5675 2431
rect 5917 2397 5951 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 8033 2397 8067 2431
rect 9229 2397 9263 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 11069 2397 11103 2431
rect 11345 2397 11379 2431
rect 3157 2329 3191 2363
rect 6561 2329 6595 2363
rect 9321 2261 9355 2295
<< metal1 >>
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 8662 12628 8668 12640
rect 7800 12600 8668 12628
rect 7800 12588 7806 12600
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 1104 12538 11868 12560
rect 1104 12486 2295 12538
rect 2347 12486 2359 12538
rect 2411 12486 2423 12538
rect 2475 12486 2487 12538
rect 2539 12486 2551 12538
rect 2603 12486 4986 12538
rect 5038 12486 5050 12538
rect 5102 12486 5114 12538
rect 5166 12486 5178 12538
rect 5230 12486 5242 12538
rect 5294 12486 7677 12538
rect 7729 12486 7741 12538
rect 7793 12486 7805 12538
rect 7857 12486 7869 12538
rect 7921 12486 7933 12538
rect 7985 12486 10368 12538
rect 10420 12486 10432 12538
rect 10484 12486 10496 12538
rect 10548 12486 10560 12538
rect 10612 12486 10624 12538
rect 10676 12486 11868 12538
rect 1104 12464 11868 12486
rect 1486 12384 1492 12436
rect 1544 12384 1550 12436
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3936 12396 4077 12424
rect 3936 12384 3942 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 5592 12396 8493 12424
rect 5592 12384 5598 12396
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 12894 12424 12900 12436
rect 10275 12396 12900 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 2501 12359 2559 12365
rect 2501 12325 2513 12359
rect 2547 12356 2559 12359
rect 4890 12356 4896 12368
rect 2547 12328 4896 12356
rect 2547 12325 2559 12328
rect 2501 12319 2559 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 7558 12316 7564 12368
rect 7616 12356 7622 12368
rect 7745 12359 7803 12365
rect 7745 12356 7757 12359
rect 7616 12328 7757 12356
rect 7616 12316 7622 12328
rect 7745 12325 7757 12328
rect 7791 12325 7803 12359
rect 8389 12359 8447 12365
rect 7745 12319 7803 12325
rect 7944 12328 8248 12356
rect 14 12248 20 12300
rect 72 12288 78 12300
rect 72 12260 2360 12288
rect 72 12248 78 12260
rect 1026 12180 1032 12232
rect 1084 12220 1090 12232
rect 2332 12229 2360 12260
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 7834 12288 7840 12300
rect 4120 12260 7840 12288
rect 4120 12248 4126 12260
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1084 12192 2053 12220
rect 1084 12180 1090 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 3804 12192 4200 12220
rect 1762 12112 1768 12164
rect 1820 12112 1826 12164
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 3804 12152 3832 12192
rect 2271 12124 3832 12152
rect 4172 12152 4200 12192
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 4304 12192 4353 12220
rect 4304 12180 4310 12192
rect 4341 12189 4353 12192
rect 4387 12220 4399 12223
rect 5350 12220 5356 12232
rect 4387 12192 5356 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 6546 12180 6552 12232
rect 6604 12180 6610 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7469 12223 7527 12229
rect 7469 12220 7481 12223
rect 7340 12192 7481 12220
rect 7340 12180 7346 12192
rect 7469 12189 7481 12192
rect 7515 12220 7527 12223
rect 7944 12220 7972 12328
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8220 12288 8248 12328
rect 8389 12325 8401 12359
rect 8435 12356 8447 12359
rect 9766 12356 9772 12368
rect 8435 12328 9772 12356
rect 8435 12325 8447 12328
rect 8389 12319 8447 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 8076 12260 8156 12288
rect 8220 12260 8308 12288
rect 8076 12248 8082 12260
rect 8128 12229 8156 12260
rect 7515 12192 7972 12220
rect 8113 12223 8171 12229
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8280 12220 8308 12260
rect 8280 12192 8524 12220
rect 8113 12183 8171 12189
rect 5629 12155 5687 12161
rect 4172 12124 4660 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 4632 12084 4660 12124
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 6270 12152 6276 12164
rect 5675 12124 6276 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 7944 12124 8401 12152
rect 7944 12096 7972 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 8496 12152 8524 12192
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9646 12192 10180 12220
rect 9646 12152 9674 12192
rect 8496 12124 9674 12152
rect 9953 12155 10011 12161
rect 8389 12115 8447 12121
rect 9953 12121 9965 12155
rect 9999 12152 10011 12155
rect 10042 12152 10048 12164
rect 9999 12124 10048 12152
rect 9999 12121 10011 12124
rect 9953 12115 10011 12121
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10152 12152 10180 12192
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10284 12192 10609 12220
rect 10284 12180 10290 12192
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 10870 12152 10876 12164
rect 10152 12124 10876 12152
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 6546 12084 6552 12096
rect 4632 12056 6552 12084
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 7926 12044 7932 12096
rect 7984 12044 7990 12096
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12084 8263 12087
rect 8294 12084 8300 12096
rect 8251 12056 8300 12084
rect 8251 12053 8263 12056
rect 8205 12047 8263 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9309 12087 9367 12093
rect 9309 12084 9321 12087
rect 9180 12056 9321 12084
rect 9180 12044 9186 12056
rect 9309 12053 9321 12056
rect 9355 12053 9367 12087
rect 9309 12047 9367 12053
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 9456 12056 10517 12084
rect 9456 12044 9462 12056
rect 10505 12053 10517 12056
rect 10551 12053 10563 12087
rect 10505 12047 10563 12053
rect 1104 11994 11868 12016
rect 1104 11942 2955 11994
rect 3007 11942 3019 11994
rect 3071 11942 3083 11994
rect 3135 11942 3147 11994
rect 3199 11942 3211 11994
rect 3263 11942 5646 11994
rect 5698 11942 5710 11994
rect 5762 11942 5774 11994
rect 5826 11942 5838 11994
rect 5890 11942 5902 11994
rect 5954 11942 8337 11994
rect 8389 11942 8401 11994
rect 8453 11942 8465 11994
rect 8517 11942 8529 11994
rect 8581 11942 8593 11994
rect 8645 11942 11028 11994
rect 11080 11942 11092 11994
rect 11144 11942 11156 11994
rect 11208 11942 11220 11994
rect 11272 11942 11284 11994
rect 11336 11942 11868 11994
rect 1104 11920 11868 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 1820 11852 4476 11880
rect 1820 11840 1826 11852
rect 4246 11812 4252 11824
rect 3528 11784 4252 11812
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 3528 11753 3556 11784
rect 4246 11772 4252 11784
rect 4304 11772 4310 11824
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1360 11716 1409 11744
rect 1360 11704 1366 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 4062 11704 4068 11756
rect 4120 11704 4126 11756
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 1854 11676 1860 11688
rect 1811 11648 1860 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 2740 11648 3617 11676
rect 2740 11636 2746 11648
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 3605 11639 3663 11645
rect 3712 11648 4169 11676
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 2041 11611 2099 11617
rect 2041 11608 2053 11611
rect 1728 11580 2053 11608
rect 1728 11568 1734 11580
rect 2041 11577 2053 11580
rect 2087 11577 2099 11611
rect 2041 11571 2099 11577
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 3418 11608 3424 11620
rect 3099 11580 3424 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 3510 11568 3516 11620
rect 3568 11608 3574 11620
rect 3712 11608 3740 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4448 11676 4476 11852
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 9674 11880 9680 11892
rect 4580 11852 9680 11880
rect 4580 11840 4586 11852
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 9732 11852 10333 11880
rect 9732 11840 9738 11852
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 11606 11880 11612 11892
rect 10321 11843 10379 11849
rect 10796 11852 11612 11880
rect 5534 11772 5540 11824
rect 5592 11772 5598 11824
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6512 11784 7328 11812
rect 6512 11772 6518 11784
rect 7300 11756 7328 11784
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4580 11716 4629 11744
rect 4580 11704 4586 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 4617 11707 4675 11713
rect 6012 11716 6561 11744
rect 6012 11688 6040 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 4448 11648 5856 11676
rect 4157 11639 4215 11645
rect 5828 11617 5856 11648
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 3568 11580 3740 11608
rect 5813 11611 5871 11617
rect 3568 11568 3574 11580
rect 5813 11577 5825 11611
rect 5859 11577 5871 11611
rect 5813 11571 5871 11577
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 6840 11608 6868 11707
rect 7024 11676 7052 11707
rect 7282 11704 7288 11756
rect 7340 11704 7346 11756
rect 7926 11704 7932 11756
rect 7984 11704 7990 11756
rect 8018 11704 8024 11756
rect 8076 11704 8082 11756
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8260 11716 8708 11744
rect 8260 11704 8266 11716
rect 7374 11676 7380 11688
rect 7024 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11676 7803 11679
rect 8036 11676 8064 11704
rect 8680 11685 8708 11716
rect 8864 11716 9137 11744
rect 7791 11648 8064 11676
rect 8665 11679 8723 11685
rect 7791 11645 7803 11648
rect 7745 11639 7803 11645
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 6236 11580 6868 11608
rect 6236 11568 6242 11580
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 7156 11580 8033 11608
rect 7156 11568 7162 11580
rect 8021 11577 8033 11580
rect 8067 11577 8079 11611
rect 8864 11608 8892 11716
rect 9125 11713 9137 11716
rect 9171 11744 9183 11747
rect 9858 11744 9864 11756
rect 9171 11716 9864 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10796 11753 10824 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 11333 11815 11391 11821
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 11422 11812 11428 11824
rect 11379 11784 11428 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 10520 11676 10548 11707
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10928 11716 10977 11744
rect 10928 11704 10934 11716
rect 10965 11713 10977 11716
rect 11011 11744 11023 11747
rect 11606 11744 11612 11756
rect 11011 11716 11612 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11606 11704 11612 11716
rect 11664 11704 11670 11756
rect 11514 11676 11520 11688
rect 10520 11648 11520 11676
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 8021 11571 8079 11577
rect 8680 11580 8892 11608
rect 1578 11500 1584 11552
rect 1636 11500 1642 11552
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2004 11512 2237 11540
rect 2004 11500 2010 11512
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2225 11503 2283 11509
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3329 11543 3387 11549
rect 3329 11540 3341 11543
rect 2924 11512 3341 11540
rect 2924 11500 2930 11512
rect 3329 11509 3341 11512
rect 3375 11540 3387 11543
rect 3878 11540 3884 11552
rect 3375 11512 3884 11540
rect 3375 11509 3387 11512
rect 3329 11503 3387 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 3973 11543 4031 11549
rect 3973 11509 3985 11543
rect 4019 11540 4031 11543
rect 4246 11540 4252 11552
rect 4019 11512 4252 11540
rect 4019 11509 4031 11512
rect 3973 11503 4031 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4430 11500 4436 11552
rect 4488 11500 4494 11552
rect 6362 11500 6368 11552
rect 6420 11500 6426 11552
rect 7558 11500 7564 11552
rect 7616 11500 7622 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8680 11540 8708 11580
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 8996 11580 10609 11608
rect 8996 11568 9002 11580
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 10597 11571 10655 11577
rect 7892 11512 8708 11540
rect 7892 11500 7898 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8812 11512 9045 11540
rect 8812 11500 8818 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9398 11540 9404 11552
rect 9079 11512 9404 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 1104 11450 11868 11472
rect 1104 11398 2295 11450
rect 2347 11398 2359 11450
rect 2411 11398 2423 11450
rect 2475 11398 2487 11450
rect 2539 11398 2551 11450
rect 2603 11398 4986 11450
rect 5038 11398 5050 11450
rect 5102 11398 5114 11450
rect 5166 11398 5178 11450
rect 5230 11398 5242 11450
rect 5294 11398 7677 11450
rect 7729 11398 7741 11450
rect 7793 11398 7805 11450
rect 7857 11398 7869 11450
rect 7921 11398 7933 11450
rect 7985 11398 10368 11450
rect 10420 11398 10432 11450
rect 10484 11398 10496 11450
rect 10548 11398 10560 11450
rect 10612 11398 10624 11450
rect 10676 11398 11868 11450
rect 1104 11376 11868 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 2317 11339 2375 11345
rect 2317 11336 2329 11339
rect 2096 11308 2329 11336
rect 2096 11296 2102 11308
rect 2317 11305 2329 11308
rect 2363 11336 2375 11339
rect 2682 11336 2688 11348
rect 2363 11308 2688 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3602 11336 3608 11348
rect 3068 11308 3608 11336
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 2222 11268 2228 11280
rect 2004 11240 2228 11268
rect 2004 11228 2010 11240
rect 2222 11228 2228 11240
rect 2280 11228 2286 11280
rect 2501 11271 2559 11277
rect 2501 11237 2513 11271
rect 2547 11268 2559 11271
rect 2774 11268 2780 11280
rect 2547 11240 2780 11268
rect 2547 11237 2559 11240
rect 2501 11231 2559 11237
rect 2774 11228 2780 11240
rect 2832 11228 2838 11280
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1854 11132 1860 11144
rect 1443 11104 1860 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 2866 11132 2872 11144
rect 2823 11104 2872 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3068 11141 3096 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 7926 11336 7932 11348
rect 4479 11308 7932 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 3510 11268 3516 11280
rect 3252 11240 3516 11268
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3252 11064 3280 11240
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3467 11172 3893 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 2884 11036 3280 11064
rect 3344 11064 3372 11095
rect 3510 11092 3516 11144
rect 3568 11092 3574 11144
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3660 11104 3985 11132
rect 3660 11092 3666 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4448 11132 4476 11299
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 9784 11308 10333 11336
rect 4982 11228 4988 11280
rect 5040 11228 5046 11280
rect 5629 11271 5687 11277
rect 5629 11268 5641 11271
rect 5092 11240 5641 11268
rect 5092 11200 5120 11240
rect 5629 11237 5641 11240
rect 5675 11237 5687 11271
rect 5629 11231 5687 11237
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 9784 11268 9812 11308
rect 10321 11305 10333 11308
rect 10367 11305 10379 11339
rect 10321 11299 10379 11305
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10781 11339 10839 11345
rect 10468 11308 10732 11336
rect 10468 11296 10474 11308
rect 7524 11240 9812 11268
rect 7524 11228 7530 11240
rect 4632 11172 5120 11200
rect 4203 11104 4476 11132
rect 4525 11135 4583 11141
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 3418 11064 3424 11076
rect 3344 11036 3424 11064
rect 1857 10999 1915 11005
rect 1857 10965 1869 10999
rect 1903 10996 1915 10999
rect 1946 10996 1952 11008
rect 1903 10968 1952 10996
rect 1903 10965 1915 10968
rect 1857 10959 1915 10965
rect 1946 10956 1952 10968
rect 2004 10996 2010 11008
rect 2884 11005 2912 11036
rect 3418 11024 3424 11036
rect 3476 11024 3482 11076
rect 3786 11024 3792 11076
rect 3844 11024 3850 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4120 11036 4200 11064
rect 4120 11024 4126 11036
rect 2317 10999 2375 11005
rect 2317 10996 2329 10999
rect 2004 10968 2329 10996
rect 2004 10956 2010 10968
rect 2317 10965 2329 10968
rect 2363 10965 2375 10999
rect 2317 10959 2375 10965
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10965 2927 10999
rect 2869 10959 2927 10965
rect 3237 10999 3295 11005
rect 3237 10965 3249 10999
rect 3283 10996 3295 10999
rect 3326 10996 3332 11008
rect 3283 10968 3332 10996
rect 3283 10965 3295 10968
rect 3237 10959 3295 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 4172 10996 4200 11036
rect 4246 11024 4252 11076
rect 4304 11024 4310 11076
rect 4540 11064 4568 11095
rect 4356 11036 4568 11064
rect 4632 11064 4660 11172
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5592 11172 5733 11200
rect 5592 11160 5598 11172
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 9784 11200 9812 11240
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 10594 11268 10600 11280
rect 9999 11240 10600 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 10704 11268 10732 11308
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 10870 11336 10876 11348
rect 10827 11308 10876 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11333 11271 11391 11277
rect 11333 11268 11345 11271
rect 10704 11240 11345 11268
rect 11333 11237 11345 11240
rect 11379 11237 11391 11271
rect 11333 11231 11391 11237
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 5721 11163 5779 11169
rect 6748 11172 7696 11200
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 4764 11104 5181 11132
rect 4764 11092 4770 11104
rect 5169 11101 5181 11104
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11132 5319 11135
rect 6362 11132 6368 11144
rect 5307 11104 6368 11132
rect 5307 11101 5319 11104
rect 5261 11095 5319 11101
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 4798 11064 4804 11076
rect 4632 11036 4804 11064
rect 4356 10996 4384 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 4985 11067 5043 11073
rect 4985 11033 4997 11067
rect 5031 11064 5043 11067
rect 5534 11064 5540 11076
rect 5031 11036 5540 11064
rect 5031 11033 5043 11036
rect 4985 11027 5043 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6748 11064 6776 11172
rect 7098 11092 7104 11144
rect 7156 11092 7162 11144
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7668 11141 7696 11172
rect 9692 11172 9812 11200
rect 10060 11172 10977 11200
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7984 11104 8033 11132
rect 7984 11092 7990 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8754 11092 8760 11144
rect 8812 11092 8818 11144
rect 9692 11141 9720 11172
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 10060 11141 10088 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 6144 11036 6776 11064
rect 6825 11067 6883 11073
rect 6144 11024 6150 11036
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 6871 11036 6960 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 4172 10968 4384 10996
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 6178 10996 6184 11008
rect 4488 10968 6184 10996
rect 4488 10956 4494 10968
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 6932 10996 6960 11036
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 9493 11067 9551 11073
rect 9493 11064 9505 11067
rect 7064 11036 9505 11064
rect 7064 11024 7070 11036
rect 9493 11033 9505 11036
rect 9539 11033 9551 11067
rect 10520 11064 10548 11095
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 10980 11104 11069 11132
rect 10686 11064 10692 11076
rect 10520 11036 10692 11064
rect 9493 11027 9551 11033
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 10778 11024 10784 11076
rect 10836 11024 10842 11076
rect 7190 10996 7196 11008
rect 6932 10968 7196 10996
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 10704 10996 10732 11024
rect 10980 10996 11008 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11514 11092 11520 11144
rect 11572 11092 11578 11144
rect 10704 10968 11008 10996
rect 1104 10906 11868 10928
rect 1104 10854 2955 10906
rect 3007 10854 3019 10906
rect 3071 10854 3083 10906
rect 3135 10854 3147 10906
rect 3199 10854 3211 10906
rect 3263 10854 5646 10906
rect 5698 10854 5710 10906
rect 5762 10854 5774 10906
rect 5826 10854 5838 10906
rect 5890 10854 5902 10906
rect 5954 10854 8337 10906
rect 8389 10854 8401 10906
rect 8453 10854 8465 10906
rect 8517 10854 8529 10906
rect 8581 10854 8593 10906
rect 8645 10854 11028 10906
rect 11080 10854 11092 10906
rect 11144 10854 11156 10906
rect 11208 10854 11220 10906
rect 11272 10854 11284 10906
rect 11336 10854 11868 10906
rect 1104 10832 11868 10854
rect 2038 10752 2044 10804
rect 2096 10752 2102 10804
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2866 10792 2872 10804
rect 2455 10764 2872 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 2961 10795 3019 10801
rect 2961 10761 2973 10795
rect 3007 10792 3019 10795
rect 3786 10792 3792 10804
rect 3007 10764 3792 10792
rect 3007 10761 3019 10764
rect 2961 10755 3019 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 7374 10792 7380 10804
rect 4212 10764 7380 10792
rect 4212 10752 4218 10764
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 7926 10752 7932 10804
rect 7984 10752 7990 10804
rect 10137 10795 10195 10801
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10778 10792 10784 10804
rect 10183 10764 10784 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 2774 10684 2780 10736
rect 2832 10684 2838 10736
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 5813 10727 5871 10733
rect 5813 10724 5825 10727
rect 5040 10696 5825 10724
rect 5040 10684 5046 10696
rect 5813 10693 5825 10696
rect 5859 10724 5871 10727
rect 7285 10727 7343 10733
rect 5859 10696 6776 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1946 10616 1952 10668
rect 2004 10616 2010 10668
rect 2222 10616 2228 10668
rect 2280 10616 2286 10668
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6748 10665 6776 10696
rect 7285 10693 7297 10727
rect 7331 10724 7343 10727
rect 8202 10724 8208 10736
rect 7331 10696 8208 10724
rect 7331 10693 7343 10696
rect 7285 10687 7343 10693
rect 8202 10684 8208 10696
rect 8260 10733 8266 10736
rect 8260 10727 8323 10733
rect 8260 10693 8277 10727
rect 8311 10693 8323 10727
rect 8260 10687 8323 10693
rect 8481 10727 8539 10733
rect 8481 10693 8493 10727
rect 8527 10724 8539 10727
rect 8754 10724 8760 10736
rect 8527 10696 8760 10724
rect 8527 10693 8539 10696
rect 8481 10687 8539 10693
rect 8260 10684 8266 10687
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 6144 10628 6193 10656
rect 6144 10616 6150 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 6181 10619 6239 10625
rect 6288 10628 6653 10656
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6288 10588 6316 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 7156 10628 7573 10656
rect 7156 10616 7162 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8496 10656 8524 10687
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 9677 10727 9735 10733
rect 9677 10693 9689 10727
rect 9723 10724 9735 10727
rect 10226 10724 10232 10736
rect 9723 10696 10232 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 11241 10727 11299 10733
rect 11241 10724 11253 10727
rect 10520 10696 11253 10724
rect 8067 10628 8524 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 6052 10560 6316 10588
rect 6365 10591 6423 10597
rect 6052 10548 6058 10560
rect 6365 10557 6377 10591
rect 6411 10588 6423 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 6411 10560 7757 10588
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 2866 10480 2872 10532
rect 2924 10520 2930 10532
rect 3145 10523 3203 10529
rect 3145 10520 3157 10523
rect 2924 10492 3157 10520
rect 2924 10480 2930 10492
rect 3145 10489 3157 10492
rect 3191 10489 3203 10523
rect 3145 10483 3203 10489
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 6380 10520 6408 10551
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10008 10560 10241 10588
rect 10008 10548 10014 10560
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 6236 10492 6408 10520
rect 6457 10523 6515 10529
rect 6236 10480 6242 10492
rect 6457 10489 6469 10523
rect 6503 10520 6515 10523
rect 7006 10520 7012 10532
rect 6503 10492 7012 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1854 10452 1860 10464
rect 1627 10424 1860 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2096 10424 2973 10452
rect 2096 10412 2102 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 5994 10412 6000 10464
rect 6052 10412 6058 10464
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 6472 10452 6500 10483
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 7653 10523 7711 10529
rect 7653 10520 7665 10523
rect 7524 10492 7665 10520
rect 7524 10480 7530 10492
rect 7653 10489 7665 10492
rect 7699 10489 7711 10523
rect 7653 10483 7711 10489
rect 10042 10480 10048 10532
rect 10100 10480 10106 10532
rect 10134 10480 10140 10532
rect 10192 10520 10198 10532
rect 10520 10529 10548 10696
rect 11241 10693 11253 10696
rect 11287 10693 11299 10727
rect 11241 10687 11299 10693
rect 10870 10656 10876 10668
rect 10704 10628 10876 10656
rect 10704 10597 10732 10628
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 10192 10492 10517 10520
rect 10192 10480 10198 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10652 10492 10793 10520
rect 10652 10480 10658 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 6135 10424 6500 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6914 10412 6920 10464
rect 6972 10412 6978 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10888 10452 10916 10483
rect 10008 10424 10916 10452
rect 10008 10412 10014 10424
rect 1104 10362 11868 10384
rect 1104 10310 2295 10362
rect 2347 10310 2359 10362
rect 2411 10310 2423 10362
rect 2475 10310 2487 10362
rect 2539 10310 2551 10362
rect 2603 10310 4986 10362
rect 5038 10310 5050 10362
rect 5102 10310 5114 10362
rect 5166 10310 5178 10362
rect 5230 10310 5242 10362
rect 5294 10310 7677 10362
rect 7729 10310 7741 10362
rect 7793 10310 7805 10362
rect 7857 10310 7869 10362
rect 7921 10310 7933 10362
rect 7985 10310 10368 10362
rect 10420 10310 10432 10362
rect 10484 10310 10496 10362
rect 10548 10310 10560 10362
rect 10612 10310 10624 10362
rect 10676 10310 11868 10362
rect 1104 10288 11868 10310
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4798 10248 4804 10260
rect 4755 10220 4804 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5592 10220 5641 10248
rect 5592 10208 5598 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7340 10220 7665 10248
rect 7340 10208 7346 10220
rect 7653 10217 7665 10220
rect 7699 10248 7711 10251
rect 8294 10248 8300 10260
rect 7699 10220 8300 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10686 10248 10692 10260
rect 10551 10220 10692 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 9306 10180 9312 10192
rect 2746 10152 9312 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2746 10112 2774 10152
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 10226 10140 10232 10192
rect 10284 10180 10290 10192
rect 10321 10183 10379 10189
rect 10321 10180 10333 10183
rect 10284 10152 10333 10180
rect 10284 10140 10290 10152
rect 10321 10149 10333 10152
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 11333 10183 11391 10189
rect 11333 10149 11345 10183
rect 11379 10149 11391 10183
rect 11333 10143 11391 10149
rect 3418 10112 3424 10124
rect 1995 10084 2774 10112
rect 3068 10084 3424 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2133 10047 2191 10053
rect 2133 10044 2145 10047
rect 2096 10016 2145 10044
rect 2096 10004 2102 10016
rect 2133 10013 2145 10016
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3068 10044 3096 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4246 10072 4252 10124
rect 4304 10112 4310 10124
rect 4304 10084 5120 10112
rect 4304 10072 4310 10084
rect 2823 10016 3096 10044
rect 3145 10047 3203 10053
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3234 10044 3240 10056
rect 3191 10016 3240 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 5092 10053 5120 10084
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 11348 10112 11376 10143
rect 6696 10084 11376 10112
rect 6696 10072 6702 10084
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 3510 9936 3516 9988
rect 3568 9936 3574 9988
rect 4430 9936 4436 9988
rect 4488 9936 4494 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 4540 9908 4568 10007
rect 5442 10004 5448 10056
rect 5500 10004 5506 10056
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 7282 10044 7288 10056
rect 6052 10016 7288 10044
rect 6052 10004 6058 10016
rect 7282 10004 7288 10016
rect 7340 10044 7346 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7340 10016 7389 10044
rect 7340 10004 7346 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 5258 9936 5264 9988
rect 5316 9936 5322 9988
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 6822 9976 6828 9988
rect 5399 9948 6828 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 7685 9979 7743 9985
rect 7685 9945 7697 9979
rect 7731 9976 7743 9979
rect 8220 9976 8248 10004
rect 7731 9948 8248 9976
rect 7731 9945 7743 9948
rect 7685 9939 7743 9945
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10778 9976 10784 9988
rect 10100 9948 10784 9976
rect 10100 9936 10106 9948
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 4614 9908 4620 9920
rect 1627 9880 4620 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 7282 9908 7288 9920
rect 7239 9880 7288 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7834 9868 7840 9920
rect 7892 9868 7898 9920
rect 8018 9868 8024 9920
rect 8076 9868 8082 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 11606 9908 11612 9920
rect 10376 9880 11612 9908
rect 10376 9868 10382 9880
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 1104 9818 11868 9840
rect 1104 9766 2955 9818
rect 3007 9766 3019 9818
rect 3071 9766 3083 9818
rect 3135 9766 3147 9818
rect 3199 9766 3211 9818
rect 3263 9766 5646 9818
rect 5698 9766 5710 9818
rect 5762 9766 5774 9818
rect 5826 9766 5838 9818
rect 5890 9766 5902 9818
rect 5954 9766 8337 9818
rect 8389 9766 8401 9818
rect 8453 9766 8465 9818
rect 8517 9766 8529 9818
rect 8581 9766 8593 9818
rect 8645 9766 11028 9818
rect 11080 9766 11092 9818
rect 11144 9766 11156 9818
rect 11208 9766 11220 9818
rect 11272 9766 11284 9818
rect 11336 9766 11868 9818
rect 1104 9744 11868 9766
rect 7282 9704 7288 9716
rect 6840 9676 7288 9704
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1728 9608 3464 9636
rect 1728 9596 1734 9608
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1872 9540 2329 9568
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1872 9373 1900 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3436 9577 3464 9608
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 4154 9636 4160 9648
rect 3936 9608 4160 9636
rect 3936 9596 3942 9608
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4706 9596 4712 9648
rect 4764 9636 4770 9648
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4764 9608 4813 9636
rect 4764 9596 4770 9608
rect 4801 9605 4813 9608
rect 4847 9605 4859 9639
rect 4801 9599 4859 9605
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 5592 9608 5917 9636
rect 5592 9596 5598 9608
rect 5905 9605 5917 9608
rect 5951 9605 5963 9639
rect 6840 9636 6868 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 8018 9704 8024 9716
rect 7524 9676 8024 9704
rect 7524 9664 7530 9676
rect 8018 9664 8024 9676
rect 8076 9704 8082 9716
rect 8076 9676 8708 9704
rect 8076 9664 8082 9676
rect 8680 9636 8708 9676
rect 9214 9636 9220 9648
rect 5905 9599 5963 9605
rect 6012 9608 6868 9636
rect 6932 9608 8616 9636
rect 8680 9608 9220 9636
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2924 9540 3341 9568
rect 2924 9528 2930 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3344 9500 3372 9531
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4488 9540 4537 9568
rect 4488 9528 4494 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 3786 9500 3792 9512
rect 3344 9472 3792 9500
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4540 9500 4568 9531
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 5718 9568 5724 9580
rect 4908 9540 5724 9568
rect 4212 9472 4568 9500
rect 4212 9460 4218 9472
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 4908 9500 4936 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6012 9568 6040 9608
rect 6932 9580 6960 9608
rect 5859 9540 6040 9568
rect 6089 9571 6147 9577
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 4856 9472 4936 9500
rect 4856 9460 4862 9472
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5828 9500 5856 9531
rect 5500 9472 5856 9500
rect 6104 9500 6132 9531
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 6914 9568 6920 9580
rect 6871 9540 6920 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7466 9568 7472 9580
rect 7064 9540 7472 9568
rect 7064 9528 7070 9540
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8202 9568 8208 9580
rect 7883 9540 8208 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6104 9472 6377 9500
rect 5500 9460 5506 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 6512 9472 6745 9500
rect 6512 9460 6518 9472
rect 6733 9469 6745 9472
rect 6779 9500 6791 9503
rect 7190 9500 7196 9512
rect 6779 9472 7196 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 7576 9432 7604 9531
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 8588 9577 8616 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 8846 9568 8852 9580
rect 8619 9540 8852 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7699 9472 8125 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 9048 9500 9076 9531
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9824 9540 10149 9568
rect 9824 9528 9830 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 8812 9472 9076 9500
rect 8812 9460 8818 9472
rect 3743 9404 7604 9432
rect 7745 9435 7803 9441
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 7745 9401 7757 9435
rect 7791 9432 7803 9435
rect 7834 9432 7840 9444
rect 7791 9404 7840 9432
rect 7791 9401 7803 9404
rect 7745 9395 7803 9401
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 7944 9404 8493 9432
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1636 9336 1869 9364
rect 1636 9324 1642 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 2188 9336 2237 9364
rect 2188 9324 2194 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 3234 9364 3240 9376
rect 2455 9336 3240 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 4062 9364 4068 9376
rect 3568 9336 4068 9364
rect 3568 9324 3574 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4522 9364 4528 9376
rect 4387 9336 4528 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4522 9324 4528 9336
rect 4580 9364 4586 9376
rect 5258 9364 5264 9376
rect 4580 9336 5264 9364
rect 4580 9324 4586 9336
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5534 9324 5540 9376
rect 5592 9324 5598 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 7006 9364 7012 9376
rect 5776 9336 7012 9364
rect 5776 9324 5782 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7944 9364 7972 9404
rect 8481 9401 8493 9404
rect 8527 9432 8539 9435
rect 9030 9432 9036 9444
rect 8527 9404 9036 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 7248 9336 7972 9364
rect 7248 9324 7254 9336
rect 8018 9324 8024 9376
rect 8076 9324 8082 9376
rect 8662 9324 8668 9376
rect 8720 9324 8726 9376
rect 8941 9367 8999 9373
rect 8941 9333 8953 9367
rect 8987 9364 8999 9367
rect 9582 9364 9588 9376
rect 8987 9336 9588 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10318 9364 10324 9376
rect 10008 9336 10324 9364
rect 10008 9324 10014 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 10686 9364 10692 9376
rect 10643 9336 10692 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 1104 9274 11868 9296
rect 1104 9222 2295 9274
rect 2347 9222 2359 9274
rect 2411 9222 2423 9274
rect 2475 9222 2487 9274
rect 2539 9222 2551 9274
rect 2603 9222 4986 9274
rect 5038 9222 5050 9274
rect 5102 9222 5114 9274
rect 5166 9222 5178 9274
rect 5230 9222 5242 9274
rect 5294 9222 7677 9274
rect 7729 9222 7741 9274
rect 7793 9222 7805 9274
rect 7857 9222 7869 9274
rect 7921 9222 7933 9274
rect 7985 9222 10368 9274
rect 10420 9222 10432 9274
rect 10484 9222 10496 9274
rect 10548 9222 10560 9274
rect 10612 9222 10624 9274
rect 10676 9222 11868 9274
rect 1104 9200 11868 9222
rect 5077 9163 5135 9169
rect 5077 9129 5089 9163
rect 5123 9160 5135 9163
rect 5442 9160 5448 9172
rect 5123 9132 5448 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 8294 9160 8300 9172
rect 6788 9132 8300 9160
rect 6788 9120 6794 9132
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 9030 9120 9036 9172
rect 9088 9120 9094 9172
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 3326 9092 3332 9104
rect 2547 9064 3332 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 7926 9092 7932 9104
rect 3844 9064 7932 9092
rect 3844 9052 3850 9064
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 2188 8996 2237 9024
rect 2188 8984 2194 8996
rect 2225 8993 2237 8996
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2740 8996 2881 9024
rect 2740 8984 2746 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2777 8959 2835 8965
rect 2777 8956 2789 8959
rect 2556 8928 2789 8956
rect 2556 8916 2562 8928
rect 2777 8925 2789 8928
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 5552 8965 5580 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 8205 9095 8263 9101
rect 8205 9092 8217 9095
rect 8168 9064 8217 9092
rect 8168 9052 8174 9064
rect 8205 9061 8217 9064
rect 8251 9061 8263 9095
rect 8312 9092 8340 9120
rect 9766 9092 9772 9104
rect 8312 9064 9772 9092
rect 8205 9055 8263 9061
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 9950 9052 9956 9104
rect 10008 9092 10014 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 10008 9064 10057 9092
rect 10008 9052 10014 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 8343 8996 9413 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 4120 8928 5457 8956
rect 4120 8916 4126 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 6178 8956 6184 8968
rect 5767 8928 6184 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 4614 8848 4620 8900
rect 4672 8888 4678 8900
rect 4893 8891 4951 8897
rect 4893 8888 4905 8891
rect 4672 8860 4905 8888
rect 4672 8848 4678 8860
rect 4893 8857 4905 8860
rect 4939 8857 4951 8891
rect 5460 8888 5488 8919
rect 6178 8916 6184 8928
rect 6236 8956 6242 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 6236 8928 8125 8956
rect 6236 8916 6242 8928
rect 8113 8925 8125 8928
rect 8159 8956 8171 8959
rect 8202 8956 8208 8968
rect 8159 8928 8208 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8662 8956 8668 8968
rect 8435 8928 8668 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8904 8928 8953 8956
rect 8904 8916 8910 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9950 8956 9956 8968
rect 9263 8928 9956 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10244 8956 10272 8987
rect 10686 8984 10692 9036
rect 10744 8984 10750 9036
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10244 8928 10333 8956
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10469 8959 10527 8965
rect 10469 8925 10481 8959
rect 10515 8956 10527 8959
rect 10704 8956 10732 8984
rect 10515 8928 10732 8956
rect 10786 8959 10844 8965
rect 10515 8925 10527 8928
rect 10469 8919 10527 8925
rect 10786 8925 10798 8959
rect 10832 8925 10844 8959
rect 10786 8919 10844 8925
rect 9582 8888 9588 8900
rect 5460 8860 9588 8888
rect 4893 8851 4951 8857
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 10686 8848 10692 8900
rect 10744 8848 10750 8900
rect 10796 8832 10824 8919
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 3418 8820 3424 8832
rect 1820 8792 3424 8820
rect 1820 8780 1826 8792
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 5093 8823 5151 8829
rect 5093 8820 5105 8823
rect 4856 8792 5105 8820
rect 4856 8780 4862 8792
rect 5093 8789 5105 8792
rect 5139 8789 5151 8823
rect 5093 8783 5151 8789
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 6178 8820 6184 8832
rect 5408 8792 6184 8820
rect 5408 8780 5414 8792
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 6730 8820 6736 8832
rect 6604 8792 6736 8820
rect 6604 8780 6610 8792
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7929 8823 7987 8829
rect 7929 8789 7941 8823
rect 7975 8820 7987 8823
rect 8110 8820 8116 8832
rect 7975 8792 8116 8820
rect 7975 8789 7987 8792
rect 7929 8783 7987 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10778 8820 10784 8832
rect 9364 8792 10784 8820
rect 9364 8780 9370 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 10965 8823 11023 8829
rect 10965 8820 10977 8823
rect 10928 8792 10977 8820
rect 10928 8780 10934 8792
rect 10965 8789 10977 8792
rect 11011 8789 11023 8823
rect 10965 8783 11023 8789
rect 1104 8730 11868 8752
rect 1104 8678 2955 8730
rect 3007 8678 3019 8730
rect 3071 8678 3083 8730
rect 3135 8678 3147 8730
rect 3199 8678 3211 8730
rect 3263 8678 5646 8730
rect 5698 8678 5710 8730
rect 5762 8678 5774 8730
rect 5826 8678 5838 8730
rect 5890 8678 5902 8730
rect 5954 8678 8337 8730
rect 8389 8678 8401 8730
rect 8453 8678 8465 8730
rect 8517 8678 8529 8730
rect 8581 8678 8593 8730
rect 8645 8678 11028 8730
rect 11080 8678 11092 8730
rect 11144 8678 11156 8730
rect 11208 8678 11220 8730
rect 11272 8678 11284 8730
rect 11336 8678 11868 8730
rect 1104 8656 11868 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1670 8616 1676 8628
rect 1627 8588 1676 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2188 8588 3188 8616
rect 2188 8576 2194 8588
rect 2038 8508 2044 8560
rect 2096 8548 2102 8560
rect 2317 8551 2375 8557
rect 2317 8548 2329 8551
rect 2096 8520 2329 8548
rect 2096 8508 2102 8520
rect 2317 8517 2329 8520
rect 2363 8517 2375 8551
rect 2317 8511 2375 8517
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 2685 8551 2743 8557
rect 2685 8548 2697 8551
rect 2556 8520 2697 8548
rect 2556 8508 2562 8520
rect 2685 8517 2697 8520
rect 2731 8517 2743 8551
rect 2685 8511 2743 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2130 8440 2136 8492
rect 2188 8480 2194 8492
rect 2516 8480 2544 8508
rect 2188 8452 2544 8480
rect 2593 8483 2651 8489
rect 2188 8440 2194 8452
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2608 8344 2636 8443
rect 2774 8440 2780 8492
rect 2832 8440 2838 8492
rect 3160 8489 3188 8588
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6638 8616 6644 8628
rect 6052 8588 6644 8616
rect 6052 8576 6058 8588
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8478 8616 8484 8628
rect 7984 8588 8484 8616
rect 7984 8576 7990 8588
rect 8478 8576 8484 8588
rect 8536 8616 8542 8628
rect 8754 8616 8760 8628
rect 8536 8588 8760 8616
rect 8536 8576 8542 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9214 8616 9220 8628
rect 8996 8588 9220 8616
rect 8996 8576 9002 8588
rect 9214 8576 9220 8588
rect 9272 8616 9278 8628
rect 9559 8619 9617 8625
rect 9559 8616 9571 8619
rect 9272 8588 9571 8616
rect 9272 8576 9278 8588
rect 9559 8585 9571 8588
rect 9605 8585 9617 8619
rect 9559 8579 9617 8585
rect 10321 8619 10379 8625
rect 10321 8585 10333 8619
rect 10367 8616 10379 8619
rect 10594 8616 10600 8628
rect 10367 8588 10600 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 10928 8588 11253 8616
rect 10928 8576 10934 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11241 8579 11299 8585
rect 3878 8548 3884 8560
rect 3252 8520 3884 8548
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 3252 8412 3280 8520
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4706 8548 4712 8560
rect 4540 8520 4712 8548
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 3697 8483 3755 8489
rect 3467 8452 3648 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3099 8384 3280 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3620 8412 3648 8452
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4246 8480 4252 8492
rect 3743 8452 4252 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4246 8440 4252 8452
rect 4304 8480 4310 8492
rect 4540 8489 4568 8520
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 5537 8551 5595 8557
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 6178 8548 6184 8560
rect 5583 8520 6184 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 6178 8508 6184 8520
rect 6236 8508 6242 8560
rect 6822 8548 6828 8560
rect 6656 8520 6828 8548
rect 4525 8483 4583 8489
rect 4304 8452 4476 8480
rect 4304 8440 4310 8452
rect 4154 8412 4160 8424
rect 3620 8384 4160 8412
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4448 8421 4476 8452
rect 4525 8449 4537 8483
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4672 8452 5089 8480
rect 4672 8440 4678 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5258 8440 5264 8492
rect 5316 8440 5322 8492
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 5644 8412 5672 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6104 8452 6377 8480
rect 6104 8412 6132 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6656 8489 6684 8520
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 7098 8548 7104 8560
rect 6880 8520 7104 8548
rect 6880 8508 6886 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 7340 8520 9168 8548
rect 7340 8508 7346 8520
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7006 8480 7012 8492
rect 6788 8452 7012 8480
rect 6788 8440 6794 8452
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 4479 8384 6132 8412
rect 6181 8415 6239 8421
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 7392 8412 7420 8443
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9140 8489 9168 8520
rect 9306 8508 9312 8560
rect 9364 8508 9370 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10226 8548 10232 8560
rect 9815 8520 10232 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 11057 8551 11115 8557
rect 11057 8517 11069 8551
rect 11103 8548 11115 8551
rect 11422 8548 11428 8560
rect 11103 8520 11428 8548
rect 11103 8517 11115 8520
rect 11057 8511 11115 8517
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8996 8452 9045 8480
rect 8996 8440 9002 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9398 8480 9404 8492
rect 9171 8452 9404 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 9950 8480 9956 8492
rect 9907 8452 9956 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 10100 8452 10425 8480
rect 10100 8440 10106 8452
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 11011 8452 11345 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11333 8449 11345 8452
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 6227 8384 7420 8412
rect 7653 8415 7711 8421
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 7699 8384 11100 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 2608 8316 3893 8344
rect 3881 8313 3893 8316
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 6086 8344 6092 8356
rect 5215 8316 6092 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 11072 8353 11100 8384
rect 9401 8347 9459 8353
rect 9401 8344 9413 8347
rect 9272 8316 9413 8344
rect 9272 8304 9278 8316
rect 9401 8313 9413 8316
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8313 11115 8347
rect 11057 8307 11115 8313
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 2961 8279 3019 8285
rect 2961 8276 2973 8279
rect 1544 8248 2973 8276
rect 1544 8236 1550 8248
rect 2961 8245 2973 8248
rect 3007 8245 3019 8279
rect 2961 8239 3019 8245
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 4948 8248 5733 8276
rect 4948 8236 4954 8248
rect 5721 8245 5733 8248
rect 5767 8276 5779 8279
rect 6546 8276 6552 8288
rect 5767 8248 6552 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 7190 8236 7196 8288
rect 7248 8236 7254 8288
rect 7558 8236 7564 8288
rect 7616 8236 7622 8288
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9585 8279 9643 8285
rect 9585 8276 9597 8279
rect 9548 8248 9597 8276
rect 9548 8236 9554 8248
rect 9585 8245 9597 8248
rect 9631 8245 9643 8279
rect 9585 8239 9643 8245
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9916 8248 9965 8276
rect 9916 8236 9922 8248
rect 9953 8245 9965 8248
rect 9999 8245 10011 8279
rect 9953 8239 10011 8245
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10870 8276 10876 8288
rect 10551 8248 10876 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 1104 8186 11868 8208
rect 1104 8134 2295 8186
rect 2347 8134 2359 8186
rect 2411 8134 2423 8186
rect 2475 8134 2487 8186
rect 2539 8134 2551 8186
rect 2603 8134 4986 8186
rect 5038 8134 5050 8186
rect 5102 8134 5114 8186
rect 5166 8134 5178 8186
rect 5230 8134 5242 8186
rect 5294 8134 7677 8186
rect 7729 8134 7741 8186
rect 7793 8134 7805 8186
rect 7857 8134 7869 8186
rect 7921 8134 7933 8186
rect 7985 8134 10368 8186
rect 10420 8134 10432 8186
rect 10484 8134 10496 8186
rect 10548 8134 10560 8186
rect 10612 8134 10624 8186
rect 10676 8134 11868 8186
rect 1104 8112 11868 8134
rect 1670 8032 1676 8084
rect 1728 8032 1734 8084
rect 2590 8032 2596 8084
rect 2648 8072 2654 8084
rect 2685 8075 2743 8081
rect 2685 8072 2697 8075
rect 2648 8044 2697 8072
rect 2648 8032 2654 8044
rect 2685 8041 2697 8044
rect 2731 8041 2743 8075
rect 2685 8035 2743 8041
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 4062 8072 4068 8084
rect 3936 8044 4068 8072
rect 3936 8032 3942 8044
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4614 8072 4620 8084
rect 4295 8044 4620 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 6086 8032 6092 8084
rect 6144 8032 6150 8084
rect 6196 8044 9444 8072
rect 1946 7964 1952 8016
rect 2004 8004 2010 8016
rect 2004 7976 2452 8004
rect 2004 7964 2010 7976
rect 2424 7936 2452 7976
rect 3234 7964 3240 8016
rect 3292 7964 3298 8016
rect 4706 8004 4712 8016
rect 3344 7976 4712 8004
rect 3344 7936 3372 7976
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 5261 8007 5319 8013
rect 5261 7973 5273 8007
rect 5307 8004 5319 8007
rect 5350 8004 5356 8016
rect 5307 7976 5356 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 2424 7908 3372 7936
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1544 7840 1961 7868
rect 1544 7828 1550 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2222 7877 2228 7880
rect 2189 7871 2228 7877
rect 2189 7837 2201 7871
rect 2189 7831 2228 7837
rect 2222 7828 2228 7831
rect 2280 7828 2286 7880
rect 2424 7877 2452 7908
rect 3068 7877 3096 7908
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 6196 7936 6224 8044
rect 6454 7964 6460 8016
rect 6512 7964 6518 8016
rect 7466 7964 7472 8016
rect 7524 7964 7530 8016
rect 8665 8007 8723 8013
rect 8665 7973 8677 8007
rect 8711 8004 8723 8007
rect 9030 8004 9036 8016
rect 8711 7976 9036 8004
rect 8711 7973 8723 7976
rect 8665 7967 8723 7973
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9214 7964 9220 8016
rect 9272 7964 9278 8016
rect 9306 7964 9312 8016
rect 9364 7964 9370 8016
rect 9416 8004 9444 8044
rect 9582 8032 9588 8084
rect 9640 8032 9646 8084
rect 11333 8007 11391 8013
rect 11333 8004 11345 8007
rect 9416 7976 11345 8004
rect 11333 7973 11345 7976
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 3568 7908 6224 7936
rect 6549 7939 6607 7945
rect 3568 7896 3574 7908
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2547 7871 2605 7877
rect 2547 7837 2559 7871
rect 2593 7868 2605 7871
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2593 7840 2973 7868
rect 2593 7837 2605 7840
rect 2547 7831 2605 7837
rect 2961 7837 2973 7840
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 3418 7868 3424 7880
rect 3375 7840 3424 7868
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 2314 7800 2320 7812
rect 1504 7772 2320 7800
rect 1504 7741 1532 7772
rect 2314 7760 2320 7772
rect 2372 7760 2378 7812
rect 2777 7803 2835 7809
rect 2777 7800 2789 7803
rect 2424 7772 2789 7800
rect 1489 7735 1547 7741
rect 1489 7701 1501 7735
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2424 7732 2452 7772
rect 2777 7769 2789 7772
rect 2823 7769 2835 7803
rect 2976 7800 3004 7831
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 3620 7877 3648 7908
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 6822 7936 6828 7948
rect 6595 7908 6828 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7190 7936 7196 7948
rect 7147 7908 7196 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3844 7840 3893 7868
rect 3844 7828 3850 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 3988 7800 4016 7831
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4120 7840 4537 7868
rect 4120 7828 4126 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 4982 7868 4988 7880
rect 4856 7840 4988 7868
rect 4856 7828 4862 7840
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5442 7868 5448 7880
rect 5123 7840 5448 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 6638 7868 6644 7880
rect 6319 7840 6644 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7064 7840 7481 7868
rect 7064 7828 7070 7840
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 4246 7800 4252 7812
rect 2976 7772 3556 7800
rect 3988 7772 4252 7800
rect 2777 7763 2835 7769
rect 2188 7704 2452 7732
rect 2188 7692 2194 7704
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 2866 7732 2872 7744
rect 2740 7704 2872 7732
rect 2740 7692 2746 7704
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3528 7741 3556 7772
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4948 7772 5273 7800
rect 4948 7760 4954 7772
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 5261 7763 5319 7769
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7732 3571 7735
rect 3694 7732 3700 7744
rect 3559 7704 3700 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 4212 7704 4445 7732
rect 4212 7692 4218 7704
rect 4433 7701 4445 7704
rect 4479 7732 4491 7735
rect 5994 7732 6000 7744
rect 4479 7704 6000 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7098 7732 7104 7744
rect 6972 7704 7104 7732
rect 6972 7692 6978 7704
rect 7098 7692 7104 7704
rect 7156 7732 7162 7744
rect 7576 7732 7604 7899
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8757 7939 8815 7945
rect 8352 7908 8616 7936
rect 8352 7896 8358 7908
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8404 7800 8432 7831
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8588 7868 8616 7908
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 8846 7936 8852 7948
rect 8803 7908 8852 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 8996 7908 9628 7936
rect 8996 7896 9002 7908
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8588 7840 9137 7868
rect 9125 7837 9137 7840
rect 9171 7868 9183 7871
rect 9214 7868 9220 7880
rect 9171 7840 9220 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9600 7877 9628 7908
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9416 7800 9444 7831
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 8404 7772 9076 7800
rect 9416 7772 9996 7800
rect 7156 7704 7604 7732
rect 7156 7692 7162 7704
rect 8202 7692 8208 7744
rect 8260 7692 8266 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9048 7732 9076 7772
rect 9582 7732 9588 7744
rect 9048 7704 9588 7732
rect 8941 7695 8999 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9968 7741 9996 7772
rect 9953 7735 10011 7741
rect 9953 7701 9965 7735
rect 9999 7701 10011 7735
rect 9953 7695 10011 7701
rect 1104 7642 11868 7664
rect 1104 7590 2955 7642
rect 3007 7590 3019 7642
rect 3071 7590 3083 7642
rect 3135 7590 3147 7642
rect 3199 7590 3211 7642
rect 3263 7590 5646 7642
rect 5698 7590 5710 7642
rect 5762 7590 5774 7642
rect 5826 7590 5838 7642
rect 5890 7590 5902 7642
rect 5954 7590 8337 7642
rect 8389 7590 8401 7642
rect 8453 7590 8465 7642
rect 8517 7590 8529 7642
rect 8581 7590 8593 7642
rect 8645 7590 11028 7642
rect 11080 7590 11092 7642
rect 11144 7590 11156 7642
rect 11208 7590 11220 7642
rect 11272 7590 11284 7642
rect 11336 7590 11868 7642
rect 1104 7568 11868 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2096 7500 2237 7528
rect 2096 7488 2102 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2832 7500 2881 7528
rect 2832 7488 2838 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 4246 7528 4252 7540
rect 3016 7500 4252 7528
rect 3016 7488 3022 7500
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5369 7531 5427 7537
rect 5369 7528 5381 7531
rect 5040 7500 5381 7528
rect 5040 7488 5046 7500
rect 5369 7497 5381 7500
rect 5415 7497 5427 7531
rect 5369 7491 5427 7497
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7558 7528 7564 7540
rect 7331 7500 7564 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9858 7528 9864 7540
rect 9088 7500 9864 7528
rect 9088 7488 9094 7500
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 3786 7460 3792 7472
rect 2372 7432 3188 7460
rect 2372 7420 2378 7432
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 2682 7392 2688 7404
rect 1872 7364 2688 7392
rect 1872 7336 1900 7364
rect 2682 7352 2688 7364
rect 2740 7392 2746 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2740 7364 2789 7392
rect 2740 7352 2746 7364
rect 2777 7361 2789 7364
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3160 7401 3188 7432
rect 3620 7432 3792 7460
rect 3620 7401 3648 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 4798 7460 4804 7472
rect 4396 7432 4804 7460
rect 4396 7420 4402 7432
rect 4798 7420 4804 7432
rect 4856 7460 4862 7472
rect 5169 7463 5227 7469
rect 5169 7460 5181 7463
rect 4856 7432 5181 7460
rect 4856 7420 4862 7432
rect 5169 7429 5181 7432
rect 5215 7429 5227 7463
rect 5169 7423 5227 7429
rect 5994 7420 6000 7472
rect 6052 7460 6058 7472
rect 7653 7463 7711 7469
rect 6052 7432 7604 7460
rect 6052 7420 6058 7432
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2222 7284 2228 7336
rect 2280 7324 2286 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 2280 7296 2329 7324
rect 2280 7284 2286 7296
rect 2317 7293 2329 7296
rect 2363 7324 2375 7327
rect 3068 7324 3096 7355
rect 3694 7352 3700 7404
rect 3752 7352 3758 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 6546 7392 6552 7404
rect 4028 7364 6552 7392
rect 4028 7352 4034 7364
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 7576 7401 7604 7432
rect 7653 7429 7665 7463
rect 7699 7460 7711 7463
rect 10962 7460 10968 7472
rect 7699 7432 10968 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 6696 7364 7481 7392
rect 6696 7352 6702 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 9766 7392 9772 7404
rect 7883 7364 9772 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 2363 7296 3096 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 5994 7324 6000 7336
rect 3476 7296 6000 7324
rect 3476 7284 3482 7296
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7852 7324 7880 7355
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 11238 7352 11244 7404
rect 11296 7352 11302 7404
rect 7432 7296 7880 7324
rect 7432 7284 7438 7296
rect 2133 7259 2191 7265
rect 2133 7225 2145 7259
rect 2179 7225 2191 7259
rect 4062 7256 4068 7268
rect 2133 7219 2191 7225
rect 2792 7228 4068 7256
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 2148 7188 2176 7219
rect 2792 7200 2820 7228
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 2685 7191 2743 7197
rect 2685 7188 2697 7191
rect 2148 7160 2697 7188
rect 2685 7157 2697 7160
rect 2731 7188 2743 7191
rect 2774 7188 2780 7200
rect 2731 7160 2780 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 3789 7191 3847 7197
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 3878 7188 3884 7200
rect 3835 7160 3884 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 3970 7148 3976 7200
rect 4028 7148 4034 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5442 7188 5448 7200
rect 5399 7160 5448 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 9916 7160 10977 7188
rect 9916 7148 9922 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 1104 7098 11868 7120
rect 1104 7046 2295 7098
rect 2347 7046 2359 7098
rect 2411 7046 2423 7098
rect 2475 7046 2487 7098
rect 2539 7046 2551 7098
rect 2603 7046 4986 7098
rect 5038 7046 5050 7098
rect 5102 7046 5114 7098
rect 5166 7046 5178 7098
rect 5230 7046 5242 7098
rect 5294 7046 7677 7098
rect 7729 7046 7741 7098
rect 7793 7046 7805 7098
rect 7857 7046 7869 7098
rect 7921 7046 7933 7098
rect 7985 7046 10368 7098
rect 10420 7046 10432 7098
rect 10484 7046 10496 7098
rect 10548 7046 10560 7098
rect 10612 7046 10624 7098
rect 10676 7046 11868 7098
rect 1104 7024 11868 7046
rect 3878 6944 3884 6996
rect 3936 6944 3942 6996
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 5442 6984 5448 6996
rect 4571 6956 5448 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 9217 6987 9275 6993
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9582 6984 9588 6996
rect 9263 6956 9588 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10502 6984 10508 6996
rect 9732 6956 10508 6984
rect 9732 6944 9738 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11422 6984 11428 6996
rect 11103 6956 11428 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 4430 6916 4436 6928
rect 1636 6888 4436 6916
rect 1636 6876 1642 6888
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 5169 6919 5227 6925
rect 5169 6885 5181 6919
rect 5215 6916 5227 6919
rect 5350 6916 5356 6928
rect 5215 6888 5356 6916
rect 5215 6885 5227 6888
rect 5169 6879 5227 6885
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 5537 6919 5595 6925
rect 5537 6885 5549 6919
rect 5583 6916 5595 6919
rect 6086 6916 6092 6928
rect 5583 6888 6092 6916
rect 5583 6885 5595 6888
rect 5537 6879 5595 6885
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 8680 6888 9168 6916
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 1544 6820 3893 6848
rect 1544 6808 1550 6820
rect 3881 6817 3893 6820
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4028 6820 5304 6848
rect 4028 6808 4034 6820
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 4890 6780 4896 6792
rect 4632 6752 4896 6780
rect 4338 6672 4344 6724
rect 4396 6672 4402 6724
rect 4546 6715 4604 6721
rect 4546 6681 4558 6715
rect 4592 6712 4604 6715
rect 4632 6712 4660 6752
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5276 6789 5304 6820
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5684 6820 5856 6848
rect 5684 6808 5690 6820
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5092 6712 5120 6743
rect 4592 6684 4660 6712
rect 4724 6684 5120 6712
rect 4592 6681 4604 6684
rect 4546 6675 4604 6681
rect 4154 6604 4160 6656
rect 4212 6604 4218 6656
rect 4724 6653 4752 6684
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4801 6647 4859 6653
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 5258 6644 5264 6656
rect 4847 6616 5264 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5460 6644 5488 6743
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5828 6789 5856 6820
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 8680 6848 8708 6888
rect 6604 6820 8708 6848
rect 6604 6808 6610 6820
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9140 6848 9168 6888
rect 10226 6876 10232 6928
rect 10284 6876 10290 6928
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 8812 6820 9076 6848
rect 9140 6820 9260 6848
rect 8812 6808 8818 6820
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 8938 6780 8944 6792
rect 6135 6752 8944 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9048 6789 9076 6820
rect 9232 6789 9260 6820
rect 10244 6820 11253 6848
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9306 6780 9312 6792
rect 9263 6752 9312 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9582 6780 9588 6792
rect 9456 6752 9588 6780
rect 9456 6740 9462 6752
rect 9582 6740 9588 6752
rect 9640 6780 9646 6792
rect 10244 6789 10272 6820
rect 9953 6783 10011 6789
rect 9953 6780 9965 6783
rect 9640 6752 9965 6780
rect 9640 6740 9646 6752
rect 9953 6749 9965 6752
rect 9999 6780 10011 6783
rect 10229 6783 10287 6789
rect 9999 6752 10180 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 6012 6712 6040 6740
rect 6454 6712 6460 6724
rect 6012 6684 6460 6712
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 10152 6712 10180 6752
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10888 6789 10916 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 10468 6752 10517 6780
rect 10468 6740 10474 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 11020 6752 11161 6780
rect 11020 6740 11026 6752
rect 11149 6749 11161 6752
rect 11195 6780 11207 6783
rect 11514 6780 11520 6792
rect 11195 6752 11520 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 10318 6712 10324 6724
rect 9548 6684 10088 6712
rect 10152 6684 10324 6712
rect 9548 6672 9554 6684
rect 10060 6656 10088 6684
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10689 6715 10747 6721
rect 10689 6681 10701 6715
rect 10735 6681 10747 6715
rect 10689 6675 10747 6681
rect 7006 6644 7012 6656
rect 5460 6616 7012 6644
rect 7006 6604 7012 6616
rect 7064 6644 7070 6656
rect 7650 6644 7656 6656
rect 7064 6616 7656 6644
rect 7064 6604 7070 6616
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 9401 6647 9459 6653
rect 9401 6613 9413 6647
rect 9447 6644 9459 6647
rect 9766 6644 9772 6656
rect 9447 6616 9772 6644
rect 9447 6613 9459 6616
rect 9401 6607 9459 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10042 6604 10048 6656
rect 10100 6604 10106 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10704 6644 10732 6675
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 10870 6644 10876 6656
rect 10468 6616 10876 6644
rect 10468 6604 10474 6616
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 1104 6554 11868 6576
rect 1104 6502 2955 6554
rect 3007 6502 3019 6554
rect 3071 6502 3083 6554
rect 3135 6502 3147 6554
rect 3199 6502 3211 6554
rect 3263 6502 5646 6554
rect 5698 6502 5710 6554
rect 5762 6502 5774 6554
rect 5826 6502 5838 6554
rect 5890 6502 5902 6554
rect 5954 6502 8337 6554
rect 8389 6502 8401 6554
rect 8453 6502 8465 6554
rect 8517 6502 8529 6554
rect 8581 6502 8593 6554
rect 8645 6502 11028 6554
rect 11080 6502 11092 6554
rect 11144 6502 11156 6554
rect 11208 6502 11220 6554
rect 11272 6502 11284 6554
rect 11336 6502 11868 6554
rect 1104 6480 11868 6502
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 4396 6412 4537 6440
rect 4396 6400 4402 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 4525 6403 4583 6409
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 5810 6440 5816 6452
rect 5040 6412 5816 6440
rect 5040 6400 5046 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 6104 6412 8125 6440
rect 6104 6372 6132 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10100 6412 10977 6440
rect 10100 6400 10106 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 2746 6344 6132 6372
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2746 6304 2774 6344
rect 7006 6332 7012 6384
rect 7064 6332 7070 6384
rect 7225 6375 7283 6381
rect 7225 6341 7237 6375
rect 7271 6372 7283 6375
rect 7271 6344 7420 6372
rect 7271 6341 7283 6344
rect 7225 6335 7283 6341
rect 2188 6276 2774 6304
rect 2188 6264 2194 6276
rect 4338 6264 4344 6316
rect 4396 6264 4402 6316
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4580 6276 4629 6304
rect 4580 6264 4586 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 7098 6304 7104 6316
rect 6135 6276 7104 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7392 6304 7420 6344
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 7745 6375 7803 6381
rect 7745 6372 7757 6375
rect 7524 6344 7757 6372
rect 7524 6332 7530 6344
rect 7745 6341 7757 6344
rect 7791 6341 7803 6375
rect 7745 6335 7803 6341
rect 7837 6375 7895 6381
rect 7837 6341 7849 6375
rect 7883 6372 7895 6375
rect 8220 6372 8248 6400
rect 7883 6344 8248 6372
rect 8389 6375 8447 6381
rect 7883 6341 7895 6344
rect 7837 6335 7895 6341
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 9122 6372 9128 6384
rect 8435 6344 9128 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 7392 6276 7604 6304
rect 7576 6248 7604 6276
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 5626 6236 5632 6248
rect 4764 6208 5632 6236
rect 4764 6196 4770 6208
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 7374 6236 7380 6248
rect 5767 6208 7380 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7852 6236 7880 6335
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 10413 6375 10471 6381
rect 9364 6344 10364 6372
rect 9364 6332 9370 6344
rect 8294 6313 8300 6316
rect 8292 6304 8300 6313
rect 8255 6276 8300 6304
rect 8292 6267 8300 6276
rect 8294 6264 8300 6267
rect 8352 6264 8358 6316
rect 8478 6264 8484 6316
rect 8536 6264 8542 6316
rect 8662 6304 8668 6316
rect 8623 6276 8668 6304
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 7616 6208 7880 6236
rect 8021 6239 8079 6245
rect 7616 6196 7622 6208
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8772 6236 8800 6267
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9272 6276 9505 6304
rect 9272 6264 9278 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 10336 6313 10364 6344
rect 10413 6341 10425 6375
rect 10459 6372 10471 6375
rect 11146 6372 11152 6384
rect 10459 6344 11152 6372
rect 10459 6341 10471 6344
rect 10413 6335 10471 6341
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 10594 6264 10600 6316
rect 10652 6304 10658 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10652 6276 10701 6304
rect 10652 6264 10658 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6294 10839 6307
rect 10870 6294 10876 6316
rect 10827 6273 10876 6294
rect 10781 6267 10876 6273
rect 10801 6266 10876 6267
rect 8067 6208 8800 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10801 6236 10829 6266
rect 10870 6264 10876 6266
rect 10928 6264 10934 6316
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 10468 6208 10829 6236
rect 10468 6196 10474 6208
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 5902 6168 5908 6180
rect 3568 6140 5908 6168
rect 3568 6128 3574 6140
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6089 6171 6147 6177
rect 6089 6168 6101 6171
rect 6052 6140 6101 6168
rect 6052 6128 6058 6140
rect 6089 6137 6101 6140
rect 6135 6137 6147 6171
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 6089 6131 6147 6137
rect 7116 6140 7481 6168
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 3476 6072 5089 6100
rect 3476 6060 3482 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 7116 6100 7144 6140
rect 7469 6137 7481 6140
rect 7515 6137 7527 6171
rect 7469 6131 7527 6137
rect 5500 6072 7144 6100
rect 7193 6103 7251 6109
rect 5500 6060 5506 6072
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7282 6100 7288 6112
rect 7239 6072 7288 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7374 6060 7380 6112
rect 7432 6060 7438 6112
rect 7484 6100 7512 6131
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 7708 6140 9444 6168
rect 7708 6128 7714 6140
rect 9214 6100 9220 6112
rect 7484 6072 9220 6100
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 9416 6100 9444 6140
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 9585 6171 9643 6177
rect 9585 6168 9597 6171
rect 9548 6140 9597 6168
rect 9548 6128 9554 6140
rect 9585 6137 9597 6140
rect 9631 6137 9643 6171
rect 9585 6131 9643 6137
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 10781 6171 10839 6177
rect 10781 6168 10793 6171
rect 9723 6140 10793 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10781 6137 10793 6140
rect 10827 6137 10839 6171
rect 10781 6131 10839 6137
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9416 6072 10149 6100
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 11054 6100 11060 6112
rect 10376 6072 11060 6100
rect 10376 6060 10382 6072
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 1104 6010 11868 6032
rect 1104 5958 2295 6010
rect 2347 5958 2359 6010
rect 2411 5958 2423 6010
rect 2475 5958 2487 6010
rect 2539 5958 2551 6010
rect 2603 5958 4986 6010
rect 5038 5958 5050 6010
rect 5102 5958 5114 6010
rect 5166 5958 5178 6010
rect 5230 5958 5242 6010
rect 5294 5958 7677 6010
rect 7729 5958 7741 6010
rect 7793 5958 7805 6010
rect 7857 5958 7869 6010
rect 7921 5958 7933 6010
rect 7985 5958 10368 6010
rect 10420 5958 10432 6010
rect 10484 5958 10496 6010
rect 10548 5958 10560 6010
rect 10612 5958 10624 6010
rect 10676 5958 11868 6010
rect 1104 5936 11868 5958
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 6181 5899 6239 5905
rect 6181 5896 6193 5899
rect 5408 5868 6193 5896
rect 5408 5856 5414 5868
rect 6181 5865 6193 5868
rect 6227 5865 6239 5899
rect 6181 5859 6239 5865
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9769 5899 9827 5905
rect 9769 5896 9781 5899
rect 9548 5868 9781 5896
rect 9548 5856 9554 5868
rect 9769 5865 9781 5868
rect 9815 5865 9827 5899
rect 9769 5859 9827 5865
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10042 5896 10048 5908
rect 9999 5868 10048 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10652 5868 10885 5896
rect 10652 5856 10658 5868
rect 10873 5865 10885 5868
rect 10919 5896 10931 5899
rect 11146 5896 11152 5908
rect 10919 5868 11152 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 4430 5828 4436 5840
rect 4304 5800 4436 5828
rect 4304 5788 4310 5800
rect 4430 5788 4436 5800
rect 4488 5828 4494 5840
rect 5442 5828 5448 5840
rect 4488 5800 5448 5828
rect 4488 5788 4494 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 5629 5831 5687 5837
rect 5629 5828 5641 5831
rect 5592 5800 5641 5828
rect 5592 5788 5598 5800
rect 5629 5797 5641 5800
rect 5675 5797 5687 5831
rect 10226 5828 10232 5840
rect 5629 5791 5687 5797
rect 6380 5800 10232 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1762 5760 1768 5772
rect 1443 5732 1768 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3421 5763 3479 5769
rect 3421 5760 3433 5763
rect 2740 5732 3433 5760
rect 2740 5720 2746 5732
rect 3421 5729 3433 5732
rect 3467 5729 3479 5763
rect 6380 5760 6408 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 11333 5831 11391 5837
rect 11333 5828 11345 5831
rect 10704 5800 11345 5828
rect 3421 5723 3479 5729
rect 5552 5732 6408 5760
rect 6457 5763 6515 5769
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5552 5701 5580 5732
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 7282 5760 7288 5772
rect 6503 5732 7288 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4212 5664 5457 5692
rect 4212 5652 4218 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5810 5692 5816 5704
rect 5767 5664 5816 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5810 5652 5816 5664
rect 5868 5692 5874 5704
rect 6270 5692 6276 5704
rect 5868 5664 6276 5692
rect 5868 5652 5874 5664
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6549 5695 6607 5701
rect 6411 5664 6500 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 3145 5627 3203 5633
rect 2714 5596 2774 5624
rect 2746 5556 2774 5596
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 6086 5624 6092 5636
rect 3191 5596 6092 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 5534 5556 5540 5568
rect 2746 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 5994 5556 6000 5568
rect 5951 5528 6000 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6472 5556 6500 5664
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6564 5624 6592 5655
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 7006 5692 7012 5704
rect 6748 5664 7012 5692
rect 6748 5624 6776 5664
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7116 5701 7144 5732
rect 7282 5720 7288 5732
rect 7340 5760 7346 5772
rect 7929 5763 7987 5769
rect 7340 5732 7696 5760
rect 7340 5720 7346 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5692 7251 5695
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7239 5664 7481 5692
rect 7239 5661 7251 5664
rect 7193 5655 7251 5661
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 7558 5692 7564 5704
rect 7515 5664 7564 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 6564 5596 6776 5624
rect 6822 5584 6828 5636
rect 6880 5584 6886 5636
rect 7208 5624 7236 5655
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7668 5701 7696 5732
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8202 5760 8208 5772
rect 7975 5732 8208 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8202 5720 8208 5732
rect 8260 5760 8266 5772
rect 8478 5760 8484 5772
rect 8260 5732 8484 5760
rect 8260 5720 8266 5732
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 10704 5760 10732 5800
rect 11333 5797 11345 5800
rect 11379 5797 11391 5831
rect 11333 5791 11391 5797
rect 8996 5732 10732 5760
rect 8996 5720 9002 5732
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 8294 5692 8300 5704
rect 8067 5664 8300 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8294 5652 8300 5664
rect 8352 5692 8358 5704
rect 8662 5692 8668 5704
rect 8352 5664 8668 5692
rect 8352 5652 8358 5664
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 10686 5692 10692 5704
rect 9272 5664 10692 5692
rect 9272 5652 9278 5664
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11330 5692 11336 5704
rect 10827 5664 11336 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 6932 5596 7236 5624
rect 6932 5556 6960 5596
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 9921 5627 9979 5633
rect 9921 5624 9933 5627
rect 9640 5596 9933 5624
rect 9640 5584 9646 5596
rect 9921 5593 9933 5596
rect 9967 5593 9979 5627
rect 9921 5587 9979 5593
rect 10134 5584 10140 5636
rect 10192 5624 10198 5636
rect 11606 5624 11612 5636
rect 10192 5596 11612 5624
rect 10192 5584 10198 5596
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 6472 5528 6960 5556
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7282 5556 7288 5568
rect 7064 5528 7288 5556
rect 7064 5516 7070 5528
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7374 5516 7380 5568
rect 7432 5516 7438 5568
rect 10597 5559 10655 5565
rect 10597 5525 10609 5559
rect 10643 5556 10655 5559
rect 10778 5556 10784 5568
rect 10643 5528 10784 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 1104 5466 11868 5488
rect 1104 5414 2955 5466
rect 3007 5414 3019 5466
rect 3071 5414 3083 5466
rect 3135 5414 3147 5466
rect 3199 5414 3211 5466
rect 3263 5414 5646 5466
rect 5698 5414 5710 5466
rect 5762 5414 5774 5466
rect 5826 5414 5838 5466
rect 5890 5414 5902 5466
rect 5954 5414 8337 5466
rect 8389 5414 8401 5466
rect 8453 5414 8465 5466
rect 8517 5414 8529 5466
rect 8581 5414 8593 5466
rect 8645 5414 11028 5466
rect 11080 5414 11092 5466
rect 11144 5414 11156 5466
rect 11208 5414 11220 5466
rect 11272 5414 11284 5466
rect 11336 5414 11868 5466
rect 1104 5392 11868 5414
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 2332 5324 7849 5352
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 1397 5287 1455 5293
rect 1397 5284 1409 5287
rect 992 5256 1409 5284
rect 992 5244 998 5256
rect 1397 5253 1409 5256
rect 1443 5253 1455 5287
rect 1397 5247 1455 5253
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 1946 5284 1952 5296
rect 1811 5256 1952 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 1946 5244 1952 5256
rect 2004 5244 2010 5296
rect 2332 5148 2360 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 10226 5352 10232 5364
rect 7837 5315 7895 5321
rect 8128 5324 10232 5352
rect 2682 5284 2688 5296
rect 2424 5256 2688 5284
rect 2424 5225 2452 5256
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 4614 5284 4620 5296
rect 4479 5256 4620 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 5442 5244 5448 5296
rect 5500 5284 5506 5296
rect 5721 5287 5779 5293
rect 5721 5284 5733 5287
rect 5500 5256 5733 5284
rect 5500 5244 5506 5256
rect 5721 5253 5733 5256
rect 5767 5253 5779 5287
rect 5721 5247 5779 5253
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 6914 5284 6920 5296
rect 5859 5256 6920 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 7469 5287 7527 5293
rect 7469 5284 7481 5287
rect 7248 5256 7481 5284
rect 7248 5244 7254 5256
rect 7469 5253 7481 5256
rect 7515 5253 7527 5287
rect 7469 5247 7527 5253
rect 7558 5244 7564 5296
rect 7616 5244 7622 5296
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2332 5120 2697 5148
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 3804 5080 3832 5202
rect 4632 5148 4660 5244
rect 5624 5219 5682 5225
rect 5624 5185 5636 5219
rect 5670 5216 5682 5219
rect 5994 5216 6000 5228
rect 5670 5188 5856 5216
rect 5955 5188 6000 5216
rect 5670 5185 5682 5188
rect 5624 5179 5682 5185
rect 5828 5148 5856 5188
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8128 5225 8156 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 8202 5244 8208 5296
rect 8260 5244 8266 5296
rect 9306 5284 9312 5296
rect 8404 5256 9312 5284
rect 8404 5225 8432 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7340 5188 7389 5216
rect 7340 5176 7346 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7975 5219 8033 5225
rect 7975 5216 7987 5219
rect 7377 5179 7435 5185
rect 7484 5188 7987 5216
rect 7484 5160 7512 5188
rect 7975 5185 7987 5188
rect 8021 5185 8033 5219
rect 7975 5179 8033 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8388 5219 8446 5225
rect 8388 5185 8400 5219
rect 8434 5185 8446 5219
rect 8388 5179 8446 5185
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 6546 5148 6552 5160
rect 4632 5120 5598 5148
rect 5828 5120 6552 5148
rect 5350 5080 5356 5092
rect 3804 5052 5356 5080
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 4212 4984 5457 5012
rect 4212 4972 4218 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5570 5012 5598 5120
rect 6546 5108 6552 5120
rect 6604 5148 6610 5160
rect 7466 5148 7472 5160
rect 6604 5120 7472 5148
rect 6604 5108 6610 5120
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8128 5148 8156 5179
rect 7668 5120 8156 5148
rect 8496 5148 8524 5179
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 10042 5216 10048 5228
rect 8803 5188 10048 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10284 5188 10425 5216
rect 10284 5176 10290 5188
rect 10413 5185 10425 5188
rect 10459 5216 10471 5219
rect 10502 5216 10508 5228
rect 10459 5188 10508 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11422 5216 11428 5228
rect 11379 5188 11428 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8496 5120 8677 5148
rect 7190 5040 7196 5092
rect 7248 5040 7254 5092
rect 7668 5012 7696 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 7745 5083 7803 5089
rect 7745 5049 7757 5083
rect 7791 5080 7803 5083
rect 7791 5052 8708 5080
rect 7791 5049 7803 5052
rect 7745 5043 7803 5049
rect 8680 5024 8708 5052
rect 5570 4984 7696 5012
rect 5445 4975 5503 4981
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 9732 4984 10517 5012
rect 9732 4972 9738 4984
rect 10505 4981 10517 4984
rect 10551 5012 10563 5015
rect 10962 5012 10968 5024
rect 10551 4984 10968 5012
rect 10551 4981 10563 4984
rect 10505 4975 10563 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11238 5012 11244 5024
rect 11195 4984 11244 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 1104 4922 11868 4944
rect 1104 4870 2295 4922
rect 2347 4870 2359 4922
rect 2411 4870 2423 4922
rect 2475 4870 2487 4922
rect 2539 4870 2551 4922
rect 2603 4870 4986 4922
rect 5038 4870 5050 4922
rect 5102 4870 5114 4922
rect 5166 4870 5178 4922
rect 5230 4870 5242 4922
rect 5294 4870 7677 4922
rect 7729 4870 7741 4922
rect 7793 4870 7805 4922
rect 7857 4870 7869 4922
rect 7921 4870 7933 4922
rect 7985 4870 10368 4922
rect 10420 4870 10432 4922
rect 10484 4870 10496 4922
rect 10548 4870 10560 4922
rect 10612 4870 10624 4922
rect 10676 4870 11868 4922
rect 1104 4848 11868 4870
rect 1844 4811 1902 4817
rect 1844 4777 1856 4811
rect 1890 4808 1902 4811
rect 1890 4780 4292 4808
rect 1890 4777 1902 4780
rect 1844 4771 1902 4777
rect 4264 4740 4292 4780
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 4890 4808 4896 4820
rect 4396 4780 4896 4808
rect 4396 4768 4402 4780
rect 4890 4768 4896 4780
rect 4948 4808 4954 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4948 4780 5089 4808
rect 4948 4768 4954 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 7650 4808 7656 4820
rect 5077 4771 5135 4777
rect 6104 4780 7656 4808
rect 6104 4740 6132 4780
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 9030 4808 9036 4820
rect 7760 4780 9036 4808
rect 4264 4712 6132 4740
rect 6178 4700 6184 4752
rect 6236 4700 6242 4752
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 7760 4740 7788 4780
rect 9030 4768 9036 4780
rect 9088 4808 9094 4820
rect 9490 4808 9496 4820
rect 9088 4780 9496 4808
rect 9088 4768 9094 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10042 4768 10048 4820
rect 10100 4768 10106 4820
rect 7248 4712 7788 4740
rect 7248 4700 7254 4712
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 8202 4740 8208 4752
rect 7984 4712 8208 4740
rect 7984 4700 7990 4712
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 10226 4740 10232 4752
rect 8312 4712 10232 4740
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 2590 4672 2596 4684
rect 1627 4644 2596 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 6196 4672 6224 4700
rect 5792 4644 6224 4672
rect 4614 4604 4620 4616
rect 2990 4576 4620 4604
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5792 4613 5820 4644
rect 6362 4632 6368 4684
rect 6420 4672 6426 4684
rect 8312 4672 8340 4712
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 10686 4700 10692 4752
rect 10744 4740 10750 4752
rect 10744 4712 11192 4740
rect 10744 4700 10750 4712
rect 6420 4644 8340 4672
rect 6420 4632 6426 4644
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 9732 4644 10977 4672
rect 9732 4632 9738 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 5902 4613 5908 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5408 4576 5641 4604
rect 5408 4564 5414 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5767 4607 5825 4613
rect 5767 4573 5779 4607
rect 5813 4573 5825 4607
rect 5767 4567 5825 4573
rect 5859 4607 5908 4613
rect 5859 4573 5871 4607
rect 5905 4573 5908 4607
rect 5859 4567 5908 4573
rect 5902 4564 5908 4567
rect 5960 4564 5966 4616
rect 6133 4607 6191 4613
rect 6133 4573 6145 4607
rect 6179 4573 6191 4607
rect 6133 4567 6191 4573
rect 3602 4496 3608 4548
rect 3660 4496 3666 4548
rect 3789 4539 3847 4545
rect 3789 4505 3801 4539
rect 3835 4505 3847 4539
rect 3789 4499 3847 4505
rect 1302 4428 1308 4480
rect 1360 4468 1366 4480
rect 3804 4468 3832 4499
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 5994 4539 6052 4545
rect 5994 4536 6006 4539
rect 5500 4508 6006 4536
rect 5500 4496 5506 4508
rect 5994 4505 6006 4508
rect 6040 4505 6052 4539
rect 6148 4536 6176 4567
rect 6546 4564 6552 4616
rect 6604 4564 6610 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7834 4613 7840 4616
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7432 4576 7665 4604
rect 7432 4564 7438 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 7801 4607 7840 4613
rect 7801 4573 7813 4607
rect 7801 4567 7840 4573
rect 7834 4564 7840 4567
rect 7892 4564 7898 4616
rect 8202 4613 8208 4616
rect 8159 4607 8208 4613
rect 8159 4573 8171 4607
rect 8205 4573 8208 4607
rect 8159 4567 8208 4573
rect 8202 4564 8208 4567
rect 8260 4604 8266 4616
rect 8478 4604 8484 4616
rect 8260 4576 8484 4604
rect 8260 4564 8266 4576
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4604 10195 4607
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10183 4576 10425 4604
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 10413 4573 10425 4576
rect 10459 4604 10471 4607
rect 10459 4576 10732 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 6564 4536 6592 4564
rect 6148 4508 6592 4536
rect 5994 4499 6052 4505
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7926 4536 7932 4548
rect 6972 4508 7932 4536
rect 6972 4496 6978 4508
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8021 4539 8079 4545
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 9122 4536 9128 4548
rect 8067 4508 9128 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 9122 4496 9128 4508
rect 9180 4496 9186 4548
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 10318 4536 10324 4548
rect 9272 4508 10324 4536
rect 9272 4496 9278 4508
rect 10318 4496 10324 4508
rect 10376 4536 10382 4548
rect 10376 4508 10456 4536
rect 10376 4496 10382 4508
rect 1360 4440 3832 4468
rect 1360 4428 1366 4440
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 6236 4440 6285 4468
rect 6236 4428 6242 4440
rect 6273 4437 6285 4440
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 8297 4471 8355 4477
rect 8297 4468 8309 4471
rect 6604 4440 8309 4468
rect 6604 4428 6610 4440
rect 8297 4437 8309 4440
rect 8343 4437 8355 4471
rect 8297 4431 8355 4437
rect 10134 4428 10140 4480
rect 10192 4468 10198 4480
rect 10229 4471 10287 4477
rect 10229 4468 10241 4471
rect 10192 4440 10241 4468
rect 10192 4428 10198 4440
rect 10229 4437 10241 4440
rect 10275 4437 10287 4471
rect 10428 4468 10456 4508
rect 10502 4496 10508 4548
rect 10560 4496 10566 4548
rect 10597 4539 10655 4545
rect 10597 4505 10609 4539
rect 10643 4505 10655 4539
rect 10704 4536 10732 4576
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 11054 4604 11060 4616
rect 10919 4576 11060 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11164 4613 11192 4712
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11238 4564 11244 4616
rect 11296 4564 11302 4616
rect 11256 4536 11284 4564
rect 10704 4508 11284 4536
rect 10597 4499 10655 4505
rect 10612 4468 10640 4499
rect 10428 4440 10640 4468
rect 10229 4431 10287 4437
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 11425 4471 11483 4477
rect 11425 4468 11437 4471
rect 10744 4440 11437 4468
rect 10744 4428 10750 4440
rect 11425 4437 11437 4440
rect 11471 4437 11483 4471
rect 11425 4431 11483 4437
rect 1104 4378 11868 4400
rect 1104 4326 2955 4378
rect 3007 4326 3019 4378
rect 3071 4326 3083 4378
rect 3135 4326 3147 4378
rect 3199 4326 3211 4378
rect 3263 4326 5646 4378
rect 5698 4326 5710 4378
rect 5762 4326 5774 4378
rect 5826 4326 5838 4378
rect 5890 4326 5902 4378
rect 5954 4326 8337 4378
rect 8389 4326 8401 4378
rect 8453 4326 8465 4378
rect 8517 4326 8529 4378
rect 8581 4326 8593 4378
rect 8645 4326 11028 4378
rect 11080 4326 11092 4378
rect 11144 4326 11156 4378
rect 11208 4326 11220 4378
rect 11272 4326 11284 4378
rect 11336 4326 11868 4378
rect 1104 4304 11868 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 3660 4236 5488 4264
rect 3660 4224 3666 4236
rect 2682 4196 2688 4208
rect 2424 4168 2688 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 2424 4137 2452 4168
rect 2682 4156 2688 4168
rect 2740 4156 2746 4208
rect 5460 4196 5488 4236
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5592 4236 5733 4264
rect 5592 4224 5598 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 7190 4224 7196 4276
rect 7248 4224 7254 4276
rect 7650 4224 7656 4276
rect 7708 4224 7714 4276
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 7984 4236 8064 4264
rect 7984 4224 7990 4236
rect 7098 4196 7104 4208
rect 3910 4168 5396 4196
rect 5460 4168 7104 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1688 4060 1716 4091
rect 4430 4088 4436 4140
rect 4488 4088 4494 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5368 4128 5396 4168
rect 7098 4156 7104 4168
rect 7156 4196 7162 4208
rect 7208 4196 7236 4224
rect 8036 4205 8064 4236
rect 9876 4236 10916 4264
rect 8021 4199 8079 4205
rect 7156 4168 7236 4196
rect 7484 4168 7972 4196
rect 7156 4156 7162 4168
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5368 4100 5457 4128
rect 5261 4091 5319 4097
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5583 4100 5825 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 992 4032 1716 4060
rect 992 4020 998 4032
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2188 4032 2697 4060
rect 2188 4020 2194 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 1578 3952 1584 4004
rect 1636 3952 1642 4004
rect 1854 3952 1860 4004
rect 1912 3952 1918 4004
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 4540 3924 4568 4091
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4764 4032 5181 4060
rect 4764 4020 4770 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5276 4060 5304 4091
rect 5552 4060 5580 4091
rect 5276 4032 5580 4060
rect 5828 4060 5856 4091
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6178 4128 6184 4140
rect 6135 4100 6184 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6104 4060 6132 4091
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 7484 4128 7512 4168
rect 7944 4137 7972 4168
rect 8021 4165 8033 4199
rect 8067 4165 8079 4199
rect 8021 4159 8079 4165
rect 6328 4100 7512 4128
rect 6328 4088 6334 4100
rect 5828 4032 6132 4060
rect 5169 4023 5227 4029
rect 7484 3992 7512 4100
rect 7793 4131 7851 4137
rect 7793 4097 7805 4131
rect 7839 4097 7851 4131
rect 7793 4091 7851 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 7806 4060 7834 4091
rect 8110 4088 8116 4140
rect 8168 4137 8174 4140
rect 8168 4131 8207 4137
rect 8195 4097 8207 4131
rect 8168 4091 8207 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8662 4128 8668 4140
rect 8343 4100 8668 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8168 4088 8174 4091
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9876 4128 9904 4236
rect 10778 4196 10784 4208
rect 10520 4168 10784 4196
rect 10520 4137 10548 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 9456 4100 9904 4128
rect 9953 4131 10011 4137
rect 9456 4088 9462 4100
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10505 4131 10563 4137
rect 10183 4100 10456 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 8018 4060 8024 4072
rect 7806 4032 8024 4060
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 9968 4060 9996 4091
rect 9907 4032 9996 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 10100 4032 10241 4060
rect 10100 4020 10106 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 10318 4020 10324 4072
rect 10376 4020 10382 4072
rect 10428 4060 10456 4100
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10888 4128 10916 4236
rect 11241 4131 11299 4137
rect 11241 4128 11253 4131
rect 10888 4100 11253 4128
rect 10505 4091 10563 4097
rect 11241 4097 11253 4100
rect 11287 4097 11299 4131
rect 11241 4091 11299 4097
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10428 4032 10793 4060
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 9030 3992 9036 4004
rect 7484 3964 9036 3992
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 9180 3964 10977 3992
rect 9180 3952 9186 3964
rect 2740 3896 4568 3924
rect 4709 3927 4767 3933
rect 2740 3884 2746 3896
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4798 3924 4804 3936
rect 4755 3896 4804 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 6270 3924 6276 3936
rect 5500 3896 6276 3924
rect 5500 3884 5506 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 8110 3924 8116 3936
rect 6972 3896 8116 3924
rect 6972 3884 6978 3896
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 9692 3933 9720 3964
rect 10965 3961 10977 3964
rect 11011 3992 11023 3995
rect 11422 3992 11428 4004
rect 11011 3964 11428 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3893 9735 3927
rect 9677 3887 9735 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10284 3896 10701 3924
rect 10284 3884 10290 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 1104 3834 11868 3856
rect 1104 3782 2295 3834
rect 2347 3782 2359 3834
rect 2411 3782 2423 3834
rect 2475 3782 2487 3834
rect 2539 3782 2551 3834
rect 2603 3782 4986 3834
rect 5038 3782 5050 3834
rect 5102 3782 5114 3834
rect 5166 3782 5178 3834
rect 5230 3782 5242 3834
rect 5294 3782 7677 3834
rect 7729 3782 7741 3834
rect 7793 3782 7805 3834
rect 7857 3782 7869 3834
rect 7921 3782 7933 3834
rect 7985 3782 10368 3834
rect 10420 3782 10432 3834
rect 10484 3782 10496 3834
rect 10548 3782 10560 3834
rect 10612 3782 10624 3834
rect 10676 3782 11868 3834
rect 1104 3760 11868 3782
rect 2774 3720 2780 3732
rect 2332 3692 2780 3720
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 2332 3584 2360 3692
rect 2774 3680 2780 3692
rect 2832 3720 2838 3732
rect 5442 3720 5448 3732
rect 2832 3692 5448 3720
rect 2832 3680 2838 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5555 3723 5613 3729
rect 5555 3689 5567 3723
rect 5601 3720 5613 3723
rect 6546 3720 6552 3732
rect 5601 3692 6552 3720
rect 5601 3689 5613 3692
rect 5555 3683 5613 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 8665 3723 8723 3729
rect 8665 3720 8677 3723
rect 7484 3692 8677 3720
rect 1627 3556 2360 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 3326 3544 3332 3596
rect 3384 3544 3390 3596
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 5442 3584 5448 3596
rect 3660 3556 5448 3584
rect 3660 3544 3666 3556
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5500 3556 5825 3584
rect 5500 3544 5506 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 6549 3587 6607 3593
rect 5813 3547 5871 3553
rect 5920 3556 6500 3584
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4246 3516 4252 3528
rect 3835 3488 4252 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 5920 3525 5948 3556
rect 6472 3528 6500 3556
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 7484 3584 7512 3692
rect 8665 3689 8677 3692
rect 8711 3689 8723 3723
rect 8665 3683 8723 3689
rect 9122 3680 9128 3732
rect 9180 3680 9186 3732
rect 10226 3680 10232 3732
rect 10284 3680 10290 3732
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 8754 3652 8760 3664
rect 7616 3624 8340 3652
rect 7616 3612 7622 3624
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 6595 3556 7512 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6236 3488 6377 3516
rect 6236 3476 6242 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 6454 3476 6460 3528
rect 6512 3476 6518 3528
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 6823 3519 6881 3525
rect 6823 3485 6835 3519
rect 6869 3518 6881 3519
rect 6869 3490 6960 3518
rect 6869 3485 6881 3490
rect 6823 3479 6881 3485
rect 2898 3420 3280 3448
rect 3252 3380 3280 3420
rect 4798 3408 4804 3460
rect 4856 3408 4862 3460
rect 6273 3451 6331 3457
rect 6273 3448 6285 3451
rect 5644 3420 6285 3448
rect 5644 3380 5672 3420
rect 6273 3417 6285 3420
rect 6319 3417 6331 3451
rect 6932 3448 6960 3490
rect 7098 3476 7104 3528
rect 7156 3476 7162 3528
rect 7282 3476 7288 3528
rect 7340 3476 7346 3528
rect 7484 3525 7512 3556
rect 7576 3556 7849 3584
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7300 3448 7328 3476
rect 6932 3420 7328 3448
rect 6273 3411 6331 3417
rect 7374 3408 7380 3460
rect 7432 3408 7438 3460
rect 7576 3448 7604 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 8202 3544 8208 3596
rect 8260 3544 8266 3596
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8202 3448 8208 3460
rect 7484 3420 7604 3448
rect 7668 3420 8208 3448
rect 7484 3392 7512 3420
rect 3252 3352 5672 3380
rect 5997 3383 6055 3389
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 6914 3380 6920 3392
rect 6043 3352 6920 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7009 3383 7067 3389
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7466 3380 7472 3392
rect 7055 3352 7472 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7668 3389 7696 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 8312 3448 8340 3624
rect 8496 3624 8760 3652
rect 8496 3593 8524 3624
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 9401 3655 9459 3661
rect 9401 3652 9413 3655
rect 8812 3624 9413 3652
rect 8812 3612 8818 3624
rect 9401 3621 9413 3624
rect 9447 3621 9459 3655
rect 9401 3615 9459 3621
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8996 3556 9045 3584
rect 8996 3544 9002 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3584 10471 3587
rect 10686 3584 10692 3596
rect 10459 3556 10692 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 8956 3516 8984 3544
rect 8803 3488 8984 3516
rect 9217 3519 9275 3525
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 8312 3420 8953 3448
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 8941 3411 8999 3417
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3349 7711 3383
rect 7653 3343 7711 3349
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9232 3380 9260 3479
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 8168 3352 9260 3380
rect 8168 3340 8174 3352
rect 10410 3340 10416 3392
rect 10468 3340 10474 3392
rect 1104 3290 11868 3312
rect 1104 3238 2955 3290
rect 3007 3238 3019 3290
rect 3071 3238 3083 3290
rect 3135 3238 3147 3290
rect 3199 3238 3211 3290
rect 3263 3238 5646 3290
rect 5698 3238 5710 3290
rect 5762 3238 5774 3290
rect 5826 3238 5838 3290
rect 5890 3238 5902 3290
rect 5954 3238 8337 3290
rect 8389 3238 8401 3290
rect 8453 3238 8465 3290
rect 8517 3238 8529 3290
rect 8581 3238 8593 3290
rect 8645 3238 11028 3290
rect 11080 3238 11092 3290
rect 11144 3238 11156 3290
rect 11208 3238 11220 3290
rect 11272 3238 11284 3290
rect 11336 3238 11868 3290
rect 1104 3216 11868 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 2590 3176 2596 3188
rect 1811 3148 2596 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4856 3148 4905 3176
rect 4856 3136 4862 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5408 3148 5457 3176
rect 5408 3136 5414 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6086 3176 6092 3188
rect 6043 3148 6092 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7190 3176 7196 3188
rect 6288 3148 7196 3176
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 2409 3111 2467 3117
rect 2409 3108 2421 3111
rect 1728 3080 2421 3108
rect 1728 3068 1734 3080
rect 2409 3077 2421 3080
rect 2455 3077 2467 3111
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 3726 3080 5181 3108
rect 2409 3071 2467 3077
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 6288 3108 6316 3148
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7524 3148 8064 3176
rect 7524 3136 7530 3148
rect 5169 3071 5227 3077
rect 5368 3080 6316 3108
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 5368 3049 5396 3080
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 4709 3043 4767 3049
rect 2179 3012 3004 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 14 2932 20 2984
rect 72 2972 78 2984
rect 1872 2972 1900 3003
rect 72 2944 1900 2972
rect 2976 2972 3004 3012
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4755 3012 4997 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5031 3012 5273 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 3786 2972 3792 2984
rect 2976 2944 3792 2972
rect 72 2932 78 2944
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4154 2932 4160 2984
rect 4212 2932 4218 2984
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 5166 2972 5172 2984
rect 4479 2944 5172 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 2314 2864 2320 2916
rect 2372 2864 2378 2916
rect 5276 2904 5304 3003
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5810 3040 5816 3052
rect 5675 3012 5816 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6288 3040 6316 3080
rect 6917 3111 6975 3117
rect 6917 3077 6929 3111
rect 6963 3108 6975 3111
rect 7929 3111 7987 3117
rect 7929 3108 7941 3111
rect 6963 3080 7941 3108
rect 6963 3077 6975 3080
rect 6917 3071 6975 3077
rect 7929 3077 7941 3080
rect 7975 3077 7987 3111
rect 7929 3071 7987 3077
rect 6135 3012 6316 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 5920 2972 5948 3003
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6512 3012 6653 3040
rect 6512 3000 6518 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6748 2972 6776 3003
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7650 3000 7656 3052
rect 7708 3049 7714 3052
rect 7708 3043 7759 3049
rect 7708 3009 7713 3043
rect 7747 3009 7759 3043
rect 7708 3003 7759 3009
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 7883 3012 7972 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7708 3000 7714 3003
rect 5767 2944 6776 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6178 2904 6184 2916
rect 5276 2876 6184 2904
rect 6178 2864 6184 2876
rect 6236 2864 6242 2916
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 7650 2904 7656 2916
rect 6512 2876 7656 2904
rect 6512 2864 6518 2876
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 7944 2904 7972 3012
rect 8036 2972 8064 3148
rect 8846 3136 8852 3188
rect 8904 3136 8910 3188
rect 9953 3179 10011 3185
rect 9953 3145 9965 3179
rect 9999 3176 10011 3179
rect 10042 3176 10048 3188
rect 9999 3148 10048 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11606 3176 11612 3188
rect 11195 3148 11612 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 10410 3108 10416 3120
rect 8128 3080 10416 3108
rect 8128 3049 8156 3080
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 8112 3043 8170 3049
rect 8112 3009 8124 3043
rect 8158 3009 8170 3043
rect 8112 3003 8170 3009
rect 8202 3000 8208 3052
rect 8260 3000 8266 3052
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 10778 3000 10784 3052
rect 10836 3000 10842 3052
rect 11330 3000 11336 3052
rect 11388 3000 11394 3052
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8036 2944 8309 2972
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 8110 2904 8116 2916
rect 7944 2876 8116 2904
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 1544 2808 2053 2836
rect 1544 2796 1550 2808
rect 2041 2805 2053 2808
rect 2087 2805 2099 2839
rect 2041 2799 2099 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 6696 2808 7205 2836
rect 6696 2796 6702 2808
rect 7193 2805 7205 2808
rect 7239 2805 7251 2839
rect 7193 2799 7251 2805
rect 7374 2796 7380 2848
rect 7432 2836 7438 2848
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 7432 2808 7573 2836
rect 7432 2796 7438 2808
rect 7561 2805 7573 2808
rect 7607 2836 7619 2839
rect 7926 2836 7932 2848
rect 7607 2808 7932 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 7926 2796 7932 2808
rect 7984 2836 7990 2848
rect 8404 2836 8432 2935
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9769 2907 9827 2913
rect 9769 2904 9781 2907
rect 9088 2876 9781 2904
rect 9088 2864 9094 2876
rect 9769 2873 9781 2876
rect 9815 2873 9827 2907
rect 9769 2867 9827 2873
rect 7984 2808 8432 2836
rect 7984 2796 7990 2808
rect 1104 2746 11868 2768
rect 1104 2694 2295 2746
rect 2347 2694 2359 2746
rect 2411 2694 2423 2746
rect 2475 2694 2487 2746
rect 2539 2694 2551 2746
rect 2603 2694 4986 2746
rect 5038 2694 5050 2746
rect 5102 2694 5114 2746
rect 5166 2694 5178 2746
rect 5230 2694 5242 2746
rect 5294 2694 7677 2746
rect 7729 2694 7741 2746
rect 7793 2694 7805 2746
rect 7857 2694 7869 2746
rect 7921 2694 7933 2746
rect 7985 2694 10368 2746
rect 10420 2694 10432 2746
rect 10484 2694 10496 2746
rect 10548 2694 10560 2746
rect 10612 2694 10624 2746
rect 10676 2694 11868 2746
rect 1104 2672 11868 2694
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5592 2604 6009 2632
rect 5592 2592 5598 2604
rect 5997 2601 6009 2604
rect 6043 2632 6055 2635
rect 6454 2632 6460 2644
rect 6043 2604 6460 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7524 2604 7849 2632
rect 7524 2592 7530 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10008 2604 10425 2632
rect 10008 2592 10014 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10836 2604 10885 2632
rect 10836 2592 10842 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11422 2632 11428 2644
rect 11195 2604 11428 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7190 2564 7196 2576
rect 5859 2536 7196 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 11514 2564 11520 2576
rect 10183 2536 11520 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1946 2496 1952 2508
rect 1443 2468 1952 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3602 2496 3608 2508
rect 3467 2468 3608 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 5442 2456 5448 2508
rect 5500 2456 5506 2508
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7340 2468 7481 2496
rect 7340 2456 7346 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 11422 2496 11428 2508
rect 7469 2459 7527 2465
rect 10336 2468 11428 2496
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2428 3847 2431
rect 4890 2428 4896 2440
rect 3835 2400 4896 2428
rect 3835 2397 3847 2400
rect 3789 2391 3847 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5224 2400 5641 2428
rect 5224 2388 5230 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7248 2400 7389 2428
rect 7248 2388 7254 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 10336 2437 10364 2468
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8168 2400 9229 2428
rect 8168 2388 8174 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10468 2400 10609 2428
rect 10468 2388 10474 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 11606 2428 11612 2440
rect 11379 2400 11612 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 3145 2363 3203 2369
rect 2714 2332 3096 2360
rect 3068 2292 3096 2332
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 3418 2360 3424 2372
rect 3191 2332 3424 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 3418 2320 3424 2332
rect 3476 2320 3482 2372
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6512 2332 6561 2360
rect 6512 2320 6518 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 11072 2360 11100 2391
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 12894 2360 12900 2372
rect 11072 2332 12900 2360
rect 6549 2323 6607 2329
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 4706 2292 4712 2304
rect 3068 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 1104 2202 11868 2224
rect 1104 2150 2955 2202
rect 3007 2150 3019 2202
rect 3071 2150 3083 2202
rect 3135 2150 3147 2202
rect 3199 2150 3211 2202
rect 3263 2150 5646 2202
rect 5698 2150 5710 2202
rect 5762 2150 5774 2202
rect 5826 2150 5838 2202
rect 5890 2150 5902 2202
rect 5954 2150 8337 2202
rect 8389 2150 8401 2202
rect 8453 2150 8465 2202
rect 8517 2150 8529 2202
rect 8581 2150 8593 2202
rect 8645 2150 11028 2202
rect 11080 2150 11092 2202
rect 11144 2150 11156 2202
rect 11208 2150 11220 2202
rect 11272 2150 11284 2202
rect 11336 2150 11868 2202
rect 1104 2128 11868 2150
<< via1 >>
rect 7748 12588 7800 12640
rect 8668 12588 8720 12640
rect 2295 12486 2347 12538
rect 2359 12486 2411 12538
rect 2423 12486 2475 12538
rect 2487 12486 2539 12538
rect 2551 12486 2603 12538
rect 4986 12486 5038 12538
rect 5050 12486 5102 12538
rect 5114 12486 5166 12538
rect 5178 12486 5230 12538
rect 5242 12486 5294 12538
rect 7677 12486 7729 12538
rect 7741 12486 7793 12538
rect 7805 12486 7857 12538
rect 7869 12486 7921 12538
rect 7933 12486 7985 12538
rect 10368 12486 10420 12538
rect 10432 12486 10484 12538
rect 10496 12486 10548 12538
rect 10560 12486 10612 12538
rect 10624 12486 10676 12538
rect 1492 12427 1544 12436
rect 1492 12393 1501 12427
rect 1501 12393 1535 12427
rect 1535 12393 1544 12427
rect 1492 12384 1544 12393
rect 3884 12384 3936 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 5540 12384 5592 12436
rect 12900 12384 12952 12436
rect 4896 12316 4948 12368
rect 7564 12316 7616 12368
rect 20 12248 72 12300
rect 1032 12180 1084 12232
rect 4068 12248 4120 12300
rect 7840 12248 7892 12300
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 1768 12155 1820 12164
rect 1768 12121 1777 12155
rect 1777 12121 1811 12155
rect 1811 12121 1820 12155
rect 1768 12112 1820 12121
rect 4252 12180 4304 12232
rect 5356 12180 5408 12232
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 7288 12180 7340 12232
rect 8024 12248 8076 12300
rect 9772 12316 9824 12368
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 6276 12112 6328 12164
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9036 12180 9088 12232
rect 10048 12112 10100 12164
rect 10232 12180 10284 12232
rect 10876 12112 10928 12164
rect 6552 12044 6604 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8300 12044 8352 12096
rect 9128 12044 9180 12096
rect 9404 12044 9456 12096
rect 2955 11942 3007 11994
rect 3019 11942 3071 11994
rect 3083 11942 3135 11994
rect 3147 11942 3199 11994
rect 3211 11942 3263 11994
rect 5646 11942 5698 11994
rect 5710 11942 5762 11994
rect 5774 11942 5826 11994
rect 5838 11942 5890 11994
rect 5902 11942 5954 11994
rect 8337 11942 8389 11994
rect 8401 11942 8453 11994
rect 8465 11942 8517 11994
rect 8529 11942 8581 11994
rect 8593 11942 8645 11994
rect 11028 11942 11080 11994
rect 11092 11942 11144 11994
rect 11156 11942 11208 11994
rect 11220 11942 11272 11994
rect 11284 11942 11336 11994
rect 1768 11840 1820 11892
rect 1308 11704 1360 11756
rect 4252 11772 4304 11824
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 1860 11636 1912 11688
rect 2688 11636 2740 11688
rect 1676 11568 1728 11620
rect 3424 11568 3476 11620
rect 3516 11568 3568 11620
rect 4528 11840 4580 11892
rect 9680 11840 9732 11892
rect 5540 11815 5592 11824
rect 5540 11781 5549 11815
rect 5549 11781 5583 11815
rect 5583 11781 5592 11815
rect 5540 11772 5592 11781
rect 6460 11772 6512 11824
rect 4528 11704 4580 11756
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6184 11568 6236 11620
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 7380 11636 7432 11688
rect 7104 11568 7156 11620
rect 9864 11704 9916 11756
rect 11612 11840 11664 11892
rect 11428 11772 11480 11824
rect 10876 11704 10928 11756
rect 11612 11704 11664 11756
rect 11520 11636 11572 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 1952 11500 2004 11552
rect 2872 11500 2924 11552
rect 3884 11500 3936 11552
rect 4252 11500 4304 11552
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 7840 11500 7892 11552
rect 8944 11568 8996 11620
rect 8760 11500 8812 11552
rect 9404 11500 9456 11552
rect 2295 11398 2347 11450
rect 2359 11398 2411 11450
rect 2423 11398 2475 11450
rect 2487 11398 2539 11450
rect 2551 11398 2603 11450
rect 4986 11398 5038 11450
rect 5050 11398 5102 11450
rect 5114 11398 5166 11450
rect 5178 11398 5230 11450
rect 5242 11398 5294 11450
rect 7677 11398 7729 11450
rect 7741 11398 7793 11450
rect 7805 11398 7857 11450
rect 7869 11398 7921 11450
rect 7933 11398 7985 11450
rect 10368 11398 10420 11450
rect 10432 11398 10484 11450
rect 10496 11398 10548 11450
rect 10560 11398 10612 11450
rect 10624 11398 10676 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2044 11296 2096 11348
rect 2688 11296 2740 11348
rect 1952 11271 2004 11280
rect 1952 11237 1961 11271
rect 1961 11237 1995 11271
rect 1995 11237 2004 11271
rect 1952 11228 2004 11237
rect 2228 11228 2280 11280
rect 2780 11228 2832 11280
rect 1860 11092 1912 11144
rect 2872 11092 2924 11144
rect 3608 11296 3660 11348
rect 3516 11228 3568 11280
rect 3516 11135 3568 11144
rect 3516 11101 3525 11135
rect 3525 11101 3559 11135
rect 3559 11101 3568 11135
rect 3516 11092 3568 11101
rect 3608 11092 3660 11144
rect 7932 11296 7984 11348
rect 4988 11271 5040 11280
rect 4988 11237 4997 11271
rect 4997 11237 5031 11271
rect 5031 11237 5040 11271
rect 4988 11228 5040 11237
rect 7472 11228 7524 11280
rect 10416 11296 10468 11348
rect 1952 10956 2004 11008
rect 3424 11024 3476 11076
rect 3792 11067 3844 11076
rect 3792 11033 3801 11067
rect 3801 11033 3835 11067
rect 3835 11033 3844 11067
rect 3792 11024 3844 11033
rect 4068 11024 4120 11076
rect 3332 10956 3384 11008
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 5540 11160 5592 11212
rect 10600 11228 10652 11280
rect 10876 11296 10928 11348
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 6368 11092 6420 11144
rect 4804 11067 4856 11076
rect 4804 11033 4813 11067
rect 4813 11033 4847 11067
rect 4847 11033 4856 11067
rect 4804 11024 4856 11033
rect 5540 11024 5592 11076
rect 6092 11067 6144 11076
rect 6092 11033 6101 11067
rect 6101 11033 6135 11067
rect 6135 11033 6144 11067
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7932 11092 7984 11144
rect 8760 11135 8812 11144
rect 8760 11101 8769 11135
rect 8769 11101 8803 11135
rect 8803 11101 8812 11135
rect 8760 11092 8812 11101
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 6092 11024 6144 11033
rect 4436 10956 4488 11008
rect 6184 10956 6236 11008
rect 7012 11024 7064 11076
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 10692 11024 10744 11076
rect 10784 11067 10836 11076
rect 10784 11033 10793 11067
rect 10793 11033 10827 11067
rect 10827 11033 10836 11067
rect 10784 11024 10836 11033
rect 7196 10956 7248 11008
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 2955 10854 3007 10906
rect 3019 10854 3071 10906
rect 3083 10854 3135 10906
rect 3147 10854 3199 10906
rect 3211 10854 3263 10906
rect 5646 10854 5698 10906
rect 5710 10854 5762 10906
rect 5774 10854 5826 10906
rect 5838 10854 5890 10906
rect 5902 10854 5954 10906
rect 8337 10854 8389 10906
rect 8401 10854 8453 10906
rect 8465 10854 8517 10906
rect 8529 10854 8581 10906
rect 8593 10854 8645 10906
rect 11028 10854 11080 10906
rect 11092 10854 11144 10906
rect 11156 10854 11208 10906
rect 11220 10854 11272 10906
rect 11284 10854 11336 10906
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2872 10752 2924 10804
rect 3792 10752 3844 10804
rect 4160 10752 4212 10804
rect 7380 10752 7432 10804
rect 7932 10795 7984 10804
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 10784 10752 10836 10804
rect 2780 10727 2832 10736
rect 2780 10693 2789 10727
rect 2789 10693 2823 10727
rect 2823 10693 2832 10727
rect 2780 10684 2832 10693
rect 4988 10684 5040 10736
rect 940 10616 992 10668
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 6092 10616 6144 10668
rect 8208 10684 8260 10736
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 7104 10616 7156 10668
rect 8760 10684 8812 10736
rect 10232 10684 10284 10736
rect 6000 10548 6052 10557
rect 2872 10480 2924 10532
rect 6184 10480 6236 10532
rect 9956 10548 10008 10600
rect 1860 10412 1912 10464
rect 2044 10412 2096 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 7012 10480 7064 10532
rect 7472 10480 7524 10532
rect 10048 10523 10100 10532
rect 10048 10489 10057 10523
rect 10057 10489 10091 10523
rect 10091 10489 10100 10523
rect 10048 10480 10100 10489
rect 10140 10480 10192 10532
rect 10876 10616 10928 10668
rect 10600 10480 10652 10532
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 9956 10412 10008 10464
rect 2295 10310 2347 10362
rect 2359 10310 2411 10362
rect 2423 10310 2475 10362
rect 2487 10310 2539 10362
rect 2551 10310 2603 10362
rect 4986 10310 5038 10362
rect 5050 10310 5102 10362
rect 5114 10310 5166 10362
rect 5178 10310 5230 10362
rect 5242 10310 5294 10362
rect 7677 10310 7729 10362
rect 7741 10310 7793 10362
rect 7805 10310 7857 10362
rect 7869 10310 7921 10362
rect 7933 10310 7985 10362
rect 10368 10310 10420 10362
rect 10432 10310 10484 10362
rect 10496 10310 10548 10362
rect 10560 10310 10612 10362
rect 10624 10310 10676 10362
rect 4804 10208 4856 10260
rect 5540 10208 5592 10260
rect 7288 10208 7340 10260
rect 8300 10208 8352 10260
rect 10692 10208 10744 10260
rect 9312 10140 9364 10192
rect 10232 10140 10284 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2044 10004 2096 10056
rect 3424 10072 3476 10124
rect 4252 10072 4304 10124
rect 3240 10004 3292 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 6644 10072 6696 10124
rect 3516 9979 3568 9988
rect 3516 9945 3525 9979
rect 3525 9945 3559 9979
rect 3559 9945 3568 9979
rect 3516 9936 3568 9945
rect 4436 9979 4488 9988
rect 4436 9945 4445 9979
rect 4445 9945 4479 9979
rect 4479 9945 4488 9979
rect 4436 9936 4488 9945
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 6000 10004 6052 10056
rect 7288 10004 7340 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 6828 9936 6880 9988
rect 7472 9979 7524 9988
rect 7472 9945 7481 9979
rect 7481 9945 7515 9979
rect 7515 9945 7524 9979
rect 7472 9936 7524 9945
rect 10048 9979 10100 9988
rect 10048 9945 10057 9979
rect 10057 9945 10091 9979
rect 10091 9945 10100 9979
rect 10048 9936 10100 9945
rect 10784 9936 10836 9988
rect 4620 9868 4672 9920
rect 7288 9868 7340 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 10324 9868 10376 9920
rect 11612 9868 11664 9920
rect 2955 9766 3007 9818
rect 3019 9766 3071 9818
rect 3083 9766 3135 9818
rect 3147 9766 3199 9818
rect 3211 9766 3263 9818
rect 5646 9766 5698 9818
rect 5710 9766 5762 9818
rect 5774 9766 5826 9818
rect 5838 9766 5890 9818
rect 5902 9766 5954 9818
rect 8337 9766 8389 9818
rect 8401 9766 8453 9818
rect 8465 9766 8517 9818
rect 8529 9766 8581 9818
rect 8593 9766 8645 9818
rect 11028 9766 11080 9818
rect 11092 9766 11144 9818
rect 11156 9766 11208 9818
rect 11220 9766 11272 9818
rect 11284 9766 11336 9818
rect 1676 9596 1728 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 1584 9324 1636 9376
rect 2872 9528 2924 9580
rect 3884 9596 3936 9648
rect 4160 9596 4212 9648
rect 4712 9596 4764 9648
rect 5540 9596 5592 9648
rect 7288 9664 7340 9716
rect 7472 9664 7524 9716
rect 8024 9664 8076 9716
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4436 9528 4488 9580
rect 3792 9460 3844 9512
rect 4160 9460 4212 9512
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5724 9571 5776 9580
rect 4804 9460 4856 9512
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 5448 9460 5500 9512
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6920 9528 6972 9580
rect 7012 9528 7064 9580
rect 7472 9528 7524 9580
rect 6460 9460 6512 9512
rect 7196 9460 7248 9512
rect 8208 9528 8260 9580
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 9220 9596 9272 9648
rect 8852 9528 8904 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 8760 9460 8812 9512
rect 9772 9528 9824 9580
rect 7840 9392 7892 9444
rect 2136 9324 2188 9376
rect 3240 9324 3292 9376
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 4068 9324 4120 9376
rect 4528 9324 4580 9376
rect 5264 9324 5316 9376
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 5724 9324 5776 9376
rect 7012 9324 7064 9376
rect 7196 9324 7248 9376
rect 9036 9392 9088 9444
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 9588 9324 9640 9376
rect 9956 9324 10008 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 10692 9324 10744 9376
rect 2295 9222 2347 9274
rect 2359 9222 2411 9274
rect 2423 9222 2475 9274
rect 2487 9222 2539 9274
rect 2551 9222 2603 9274
rect 4986 9222 5038 9274
rect 5050 9222 5102 9274
rect 5114 9222 5166 9274
rect 5178 9222 5230 9274
rect 5242 9222 5294 9274
rect 7677 9222 7729 9274
rect 7741 9222 7793 9274
rect 7805 9222 7857 9274
rect 7869 9222 7921 9274
rect 7933 9222 7985 9274
rect 10368 9222 10420 9274
rect 10432 9222 10484 9274
rect 10496 9222 10548 9274
rect 10560 9222 10612 9274
rect 10624 9222 10676 9274
rect 5448 9120 5500 9172
rect 6736 9120 6788 9172
rect 8300 9120 8352 9172
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 3332 9052 3384 9104
rect 3792 9052 3844 9104
rect 2136 8984 2188 9036
rect 2688 8984 2740 9036
rect 2504 8916 2556 8968
rect 4068 8916 4120 8968
rect 7932 9052 7984 9104
rect 8116 9052 8168 9104
rect 9772 9052 9824 9104
rect 9956 9052 10008 9104
rect 4620 8848 4672 8900
rect 6184 8916 6236 8968
rect 8208 8916 8260 8968
rect 8668 8916 8720 8968
rect 8852 8916 8904 8968
rect 9956 8916 10008 8968
rect 10692 8984 10744 9036
rect 9588 8848 9640 8900
rect 9772 8891 9824 8900
rect 9772 8857 9781 8891
rect 9781 8857 9815 8891
rect 9815 8857 9824 8891
rect 9772 8848 9824 8857
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 10692 8891 10744 8900
rect 10692 8857 10701 8891
rect 10701 8857 10735 8891
rect 10735 8857 10744 8891
rect 10692 8848 10744 8857
rect 1768 8780 1820 8832
rect 3424 8780 3476 8832
rect 4804 8780 4856 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 5356 8780 5408 8832
rect 6184 8780 6236 8832
rect 6552 8780 6604 8832
rect 6736 8780 6788 8832
rect 8116 8780 8168 8832
rect 9312 8780 9364 8832
rect 10784 8780 10836 8832
rect 10876 8780 10928 8832
rect 2955 8678 3007 8730
rect 3019 8678 3071 8730
rect 3083 8678 3135 8730
rect 3147 8678 3199 8730
rect 3211 8678 3263 8730
rect 5646 8678 5698 8730
rect 5710 8678 5762 8730
rect 5774 8678 5826 8730
rect 5838 8678 5890 8730
rect 5902 8678 5954 8730
rect 8337 8678 8389 8730
rect 8401 8678 8453 8730
rect 8465 8678 8517 8730
rect 8529 8678 8581 8730
rect 8593 8678 8645 8730
rect 11028 8678 11080 8730
rect 11092 8678 11144 8730
rect 11156 8678 11208 8730
rect 11220 8678 11272 8730
rect 11284 8678 11336 8730
rect 1676 8576 1728 8628
rect 2136 8576 2188 8628
rect 2044 8508 2096 8560
rect 2504 8508 2556 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2136 8440 2188 8492
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 6000 8576 6052 8628
rect 6644 8576 6696 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 8760 8576 8812 8628
rect 8944 8576 8996 8628
rect 9220 8576 9272 8628
rect 10600 8576 10652 8628
rect 10876 8576 10928 8628
rect 3884 8508 3936 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 4252 8440 4304 8492
rect 4712 8508 4764 8560
rect 6184 8508 6236 8560
rect 4160 8372 4212 8424
rect 4620 8440 4672 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6828 8508 6880 8560
rect 7104 8508 7156 8560
rect 7288 8508 7340 8560
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7012 8440 7064 8492
rect 8944 8440 8996 8492
rect 9312 8551 9364 8560
rect 9312 8517 9321 8551
rect 9321 8517 9355 8551
rect 9355 8517 9364 8551
rect 9312 8508 9364 8517
rect 10232 8508 10284 8560
rect 11428 8508 11480 8560
rect 9404 8440 9456 8492
rect 9956 8440 10008 8492
rect 10048 8440 10100 8492
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 6092 8304 6144 8356
rect 9220 8304 9272 8356
rect 1492 8236 1544 8288
rect 4896 8236 4948 8288
rect 6552 8236 6604 8288
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 7564 8279 7616 8288
rect 7564 8245 7573 8279
rect 7573 8245 7607 8279
rect 7607 8245 7616 8279
rect 7564 8236 7616 8245
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 9496 8236 9548 8288
rect 9864 8236 9916 8288
rect 10876 8236 10928 8288
rect 2295 8134 2347 8186
rect 2359 8134 2411 8186
rect 2423 8134 2475 8186
rect 2487 8134 2539 8186
rect 2551 8134 2603 8186
rect 4986 8134 5038 8186
rect 5050 8134 5102 8186
rect 5114 8134 5166 8186
rect 5178 8134 5230 8186
rect 5242 8134 5294 8186
rect 7677 8134 7729 8186
rect 7741 8134 7793 8186
rect 7805 8134 7857 8186
rect 7869 8134 7921 8186
rect 7933 8134 7985 8186
rect 10368 8134 10420 8186
rect 10432 8134 10484 8186
rect 10496 8134 10548 8186
rect 10560 8134 10612 8186
rect 10624 8134 10676 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2596 8032 2648 8084
rect 3884 8032 3936 8084
rect 4068 8075 4120 8084
rect 4068 8041 4077 8075
rect 4077 8041 4111 8075
rect 4111 8041 4120 8075
rect 4068 8032 4120 8041
rect 4620 8032 4672 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 1952 7964 2004 8016
rect 3240 8007 3292 8016
rect 3240 7973 3249 8007
rect 3249 7973 3283 8007
rect 3283 7973 3292 8007
rect 3240 7964 3292 7973
rect 4712 7964 4764 8016
rect 5356 7964 5408 8016
rect 1492 7828 1544 7880
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2228 7871 2280 7880
rect 2228 7837 2235 7871
rect 2235 7837 2280 7871
rect 2228 7828 2280 7837
rect 3516 7896 3568 7948
rect 6460 8007 6512 8016
rect 6460 7973 6469 8007
rect 6469 7973 6503 8007
rect 6503 7973 6512 8007
rect 6460 7964 6512 7973
rect 7472 8007 7524 8016
rect 7472 7973 7481 8007
rect 7481 7973 7515 8007
rect 7515 7973 7524 8007
rect 7472 7964 7524 7973
rect 9036 7964 9088 8016
rect 9220 8007 9272 8016
rect 9220 7973 9229 8007
rect 9229 7973 9263 8007
rect 9263 7973 9272 8007
rect 9220 7964 9272 7973
rect 9312 8007 9364 8016
rect 9312 7973 9321 8007
rect 9321 7973 9355 8007
rect 9355 7973 9364 8007
rect 9312 7964 9364 7973
rect 9588 8075 9640 8084
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 2320 7803 2372 7812
rect 2320 7769 2329 7803
rect 2329 7769 2363 7803
rect 2363 7769 2372 7803
rect 2320 7760 2372 7769
rect 2136 7692 2188 7744
rect 3424 7828 3476 7880
rect 6828 7896 6880 7948
rect 7196 7896 7248 7948
rect 3792 7828 3844 7880
rect 4068 7828 4120 7880
rect 4804 7828 4856 7880
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5448 7828 5500 7880
rect 6644 7828 6696 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7012 7828 7064 7880
rect 2688 7692 2740 7744
rect 2872 7692 2924 7744
rect 4252 7760 4304 7812
rect 4896 7760 4948 7812
rect 3700 7692 3752 7744
rect 4160 7692 4212 7744
rect 6000 7692 6052 7744
rect 6920 7692 6972 7744
rect 7104 7692 7156 7744
rect 8300 7896 8352 7948
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8852 7896 8904 7948
rect 8944 7896 8996 7948
rect 9220 7828 9272 7880
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8668 7692 8720 7744
rect 9588 7692 9640 7744
rect 2955 7590 3007 7642
rect 3019 7590 3071 7642
rect 3083 7590 3135 7642
rect 3147 7590 3199 7642
rect 3211 7590 3263 7642
rect 5646 7590 5698 7642
rect 5710 7590 5762 7642
rect 5774 7590 5826 7642
rect 5838 7590 5890 7642
rect 5902 7590 5954 7642
rect 8337 7590 8389 7642
rect 8401 7590 8453 7642
rect 8465 7590 8517 7642
rect 8529 7590 8581 7642
rect 8593 7590 8645 7642
rect 11028 7590 11080 7642
rect 11092 7590 11144 7642
rect 11156 7590 11208 7642
rect 11220 7590 11272 7642
rect 11284 7590 11336 7642
rect 2044 7488 2096 7540
rect 2780 7488 2832 7540
rect 2964 7488 3016 7540
rect 4252 7488 4304 7540
rect 4988 7488 5040 7540
rect 7564 7488 7616 7540
rect 9036 7488 9088 7540
rect 9864 7488 9916 7540
rect 2320 7420 2372 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2688 7352 2740 7404
rect 2964 7352 3016 7404
rect 3792 7420 3844 7472
rect 4344 7420 4396 7472
rect 4804 7420 4856 7472
rect 6000 7420 6052 7472
rect 1860 7284 1912 7336
rect 2228 7284 2280 7336
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 3976 7352 4028 7404
rect 6552 7352 6604 7404
rect 6644 7352 6696 7404
rect 10968 7420 11020 7472
rect 3424 7284 3476 7336
rect 6000 7284 6052 7336
rect 7380 7284 7432 7336
rect 9772 7352 9824 7404
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 4068 7216 4120 7268
rect 2780 7148 2832 7200
rect 3884 7148 3936 7200
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 5448 7148 5500 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 9864 7148 9916 7200
rect 2295 7046 2347 7098
rect 2359 7046 2411 7098
rect 2423 7046 2475 7098
rect 2487 7046 2539 7098
rect 2551 7046 2603 7098
rect 4986 7046 5038 7098
rect 5050 7046 5102 7098
rect 5114 7046 5166 7098
rect 5178 7046 5230 7098
rect 5242 7046 5294 7098
rect 7677 7046 7729 7098
rect 7741 7046 7793 7098
rect 7805 7046 7857 7098
rect 7869 7046 7921 7098
rect 7933 7046 7985 7098
rect 10368 7046 10420 7098
rect 10432 7046 10484 7098
rect 10496 7046 10548 7098
rect 10560 7046 10612 7098
rect 10624 7046 10676 7098
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 5448 6944 5500 6996
rect 9588 6944 9640 6996
rect 9680 6944 9732 6996
rect 10508 6944 10560 6996
rect 11428 6944 11480 6996
rect 1584 6876 1636 6928
rect 4436 6876 4488 6928
rect 5356 6876 5408 6928
rect 6092 6876 6144 6928
rect 1492 6808 1544 6860
rect 3976 6808 4028 6860
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 4896 6740 4948 6792
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5632 6808 5684 6860
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 5264 6604 5316 6656
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6552 6808 6604 6860
rect 8760 6808 8812 6860
rect 10232 6919 10284 6928
rect 10232 6885 10241 6919
rect 10241 6885 10275 6919
rect 10275 6885 10284 6919
rect 10232 6876 10284 6885
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 8944 6740 8996 6792
rect 9312 6740 9364 6792
rect 9404 6740 9456 6792
rect 9588 6740 9640 6792
rect 6460 6672 6512 6724
rect 9496 6672 9548 6724
rect 10416 6740 10468 6792
rect 10968 6740 11020 6792
rect 11520 6740 11572 6792
rect 10324 6672 10376 6724
rect 7012 6604 7064 6656
rect 7656 6604 7708 6656
rect 9772 6604 9824 6656
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 10416 6604 10468 6656
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 10876 6604 10928 6656
rect 2955 6502 3007 6554
rect 3019 6502 3071 6554
rect 3083 6502 3135 6554
rect 3147 6502 3199 6554
rect 3211 6502 3263 6554
rect 5646 6502 5698 6554
rect 5710 6502 5762 6554
rect 5774 6502 5826 6554
rect 5838 6502 5890 6554
rect 5902 6502 5954 6554
rect 8337 6502 8389 6554
rect 8401 6502 8453 6554
rect 8465 6502 8517 6554
rect 8529 6502 8581 6554
rect 8593 6502 8645 6554
rect 11028 6502 11080 6554
rect 11092 6502 11144 6554
rect 11156 6502 11208 6554
rect 11220 6502 11272 6554
rect 11284 6502 11336 6554
rect 4344 6400 4396 6452
rect 4988 6400 5040 6452
rect 5816 6400 5868 6452
rect 8208 6400 8260 6452
rect 10048 6400 10100 6452
rect 2136 6264 2188 6316
rect 7012 6375 7064 6384
rect 7012 6341 7021 6375
rect 7021 6341 7055 6375
rect 7055 6341 7064 6375
rect 7012 6332 7064 6341
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4528 6264 4580 6316
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 7104 6264 7156 6316
rect 7472 6332 7524 6384
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 4712 6196 4764 6248
rect 5632 6239 5684 6248
rect 5632 6205 5641 6239
rect 5641 6205 5675 6239
rect 5675 6205 5684 6239
rect 5632 6196 5684 6205
rect 7380 6196 7432 6248
rect 7564 6196 7616 6248
rect 9128 6332 9180 6384
rect 9312 6332 9364 6384
rect 8300 6307 8352 6316
rect 8300 6273 8304 6307
rect 8304 6273 8338 6307
rect 8338 6273 8352 6307
rect 8300 6264 8352 6273
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 8668 6307 8720 6316
rect 8668 6273 8676 6307
rect 8676 6273 8710 6307
rect 8710 6273 8720 6307
rect 8668 6264 8720 6273
rect 9220 6264 9272 6316
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 11152 6332 11204 6384
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 10600 6264 10652 6316
rect 10416 6196 10468 6248
rect 10876 6264 10928 6316
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 3516 6128 3568 6180
rect 5908 6128 5960 6180
rect 6000 6128 6052 6180
rect 3424 6060 3476 6112
rect 5448 6060 5500 6112
rect 7288 6060 7340 6112
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 7656 6128 7708 6180
rect 9220 6060 9272 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 9496 6128 9548 6180
rect 10324 6060 10376 6112
rect 11060 6060 11112 6112
rect 2295 5958 2347 6010
rect 2359 5958 2411 6010
rect 2423 5958 2475 6010
rect 2487 5958 2539 6010
rect 2551 5958 2603 6010
rect 4986 5958 5038 6010
rect 5050 5958 5102 6010
rect 5114 5958 5166 6010
rect 5178 5958 5230 6010
rect 5242 5958 5294 6010
rect 7677 5958 7729 6010
rect 7741 5958 7793 6010
rect 7805 5958 7857 6010
rect 7869 5958 7921 6010
rect 7933 5958 7985 6010
rect 10368 5958 10420 6010
rect 10432 5958 10484 6010
rect 10496 5958 10548 6010
rect 10560 5958 10612 6010
rect 10624 5958 10676 6010
rect 5356 5856 5408 5908
rect 9496 5856 9548 5908
rect 10048 5856 10100 5908
rect 10600 5856 10652 5908
rect 11152 5856 11204 5908
rect 4252 5788 4304 5840
rect 4436 5788 4488 5840
rect 5448 5788 5500 5840
rect 5540 5788 5592 5840
rect 1768 5720 1820 5772
rect 2688 5720 2740 5772
rect 10232 5788 10284 5840
rect 4160 5652 4212 5704
rect 5816 5652 5868 5704
rect 6276 5652 6328 5704
rect 6092 5584 6144 5636
rect 5540 5516 5592 5568
rect 6000 5516 6052 5568
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 7012 5652 7064 5704
rect 7288 5720 7340 5772
rect 6828 5627 6880 5636
rect 6828 5593 6837 5627
rect 6837 5593 6871 5627
rect 6871 5593 6880 5627
rect 6828 5584 6880 5593
rect 7564 5652 7616 5704
rect 8208 5720 8260 5772
rect 8484 5720 8536 5772
rect 8944 5720 8996 5772
rect 8300 5652 8352 5704
rect 8668 5652 8720 5704
rect 9220 5652 9272 5704
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 11336 5652 11388 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 9588 5584 9640 5636
rect 10140 5627 10192 5636
rect 10140 5593 10149 5627
rect 10149 5593 10183 5627
rect 10183 5593 10192 5627
rect 10140 5584 10192 5593
rect 11612 5584 11664 5636
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 7288 5516 7340 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 10784 5516 10836 5568
rect 2955 5414 3007 5466
rect 3019 5414 3071 5466
rect 3083 5414 3135 5466
rect 3147 5414 3199 5466
rect 3211 5414 3263 5466
rect 5646 5414 5698 5466
rect 5710 5414 5762 5466
rect 5774 5414 5826 5466
rect 5838 5414 5890 5466
rect 5902 5414 5954 5466
rect 8337 5414 8389 5466
rect 8401 5414 8453 5466
rect 8465 5414 8517 5466
rect 8529 5414 8581 5466
rect 8593 5414 8645 5466
rect 11028 5414 11080 5466
rect 11092 5414 11144 5466
rect 11156 5414 11208 5466
rect 11220 5414 11272 5466
rect 11284 5414 11336 5466
rect 940 5244 992 5296
rect 1952 5244 2004 5296
rect 2688 5244 2740 5296
rect 4620 5244 4672 5296
rect 5448 5244 5500 5296
rect 6920 5244 6972 5296
rect 7196 5244 7248 5296
rect 7564 5287 7616 5296
rect 7564 5253 7573 5287
rect 7573 5253 7607 5287
rect 7607 5253 7616 5287
rect 7564 5244 7616 5253
rect 6000 5219 6052 5228
rect 6000 5185 6008 5219
rect 6008 5185 6042 5219
rect 6042 5185 6052 5219
rect 6000 5176 6052 5185
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 7288 5176 7340 5228
rect 10232 5312 10284 5364
rect 8208 5287 8260 5296
rect 8208 5253 8217 5287
rect 8217 5253 8251 5287
rect 8251 5253 8260 5287
rect 8208 5244 8260 5253
rect 9312 5244 9364 5296
rect 5356 5040 5408 5092
rect 4160 4972 4212 5024
rect 6552 5108 6604 5160
rect 7472 5108 7524 5160
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 10048 5176 10100 5228
rect 10232 5176 10284 5228
rect 10508 5176 10560 5228
rect 11428 5176 11480 5228
rect 7196 5083 7248 5092
rect 7196 5049 7205 5083
rect 7205 5049 7239 5083
rect 7239 5049 7248 5083
rect 7196 5040 7248 5049
rect 8668 4972 8720 5024
rect 9680 4972 9732 5024
rect 10968 4972 11020 5024
rect 11244 4972 11296 5024
rect 2295 4870 2347 4922
rect 2359 4870 2411 4922
rect 2423 4870 2475 4922
rect 2487 4870 2539 4922
rect 2551 4870 2603 4922
rect 4986 4870 5038 4922
rect 5050 4870 5102 4922
rect 5114 4870 5166 4922
rect 5178 4870 5230 4922
rect 5242 4870 5294 4922
rect 7677 4870 7729 4922
rect 7741 4870 7793 4922
rect 7805 4870 7857 4922
rect 7869 4870 7921 4922
rect 7933 4870 7985 4922
rect 10368 4870 10420 4922
rect 10432 4870 10484 4922
rect 10496 4870 10548 4922
rect 10560 4870 10612 4922
rect 10624 4870 10676 4922
rect 4344 4768 4396 4820
rect 4896 4768 4948 4820
rect 7656 4768 7708 4820
rect 6184 4700 6236 4752
rect 7196 4700 7248 4752
rect 9036 4768 9088 4820
rect 9496 4768 9548 4820
rect 10048 4811 10100 4820
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 7932 4700 7984 4752
rect 8208 4700 8260 4752
rect 2596 4632 2648 4684
rect 4620 4564 4672 4616
rect 5356 4564 5408 4616
rect 6368 4632 6420 4684
rect 10232 4700 10284 4752
rect 10692 4700 10744 4752
rect 9680 4632 9732 4684
rect 5908 4564 5960 4616
rect 3608 4539 3660 4548
rect 3608 4505 3617 4539
rect 3617 4505 3651 4539
rect 3651 4505 3660 4539
rect 3608 4496 3660 4505
rect 1308 4428 1360 4480
rect 5448 4496 5500 4548
rect 6552 4564 6604 4616
rect 7380 4564 7432 4616
rect 7840 4607 7892 4616
rect 7840 4573 7847 4607
rect 7847 4573 7892 4607
rect 7840 4564 7892 4573
rect 8208 4564 8260 4616
rect 8484 4564 8536 4616
rect 6920 4496 6972 4548
rect 7932 4539 7984 4548
rect 7932 4505 7941 4539
rect 7941 4505 7975 4539
rect 7975 4505 7984 4539
rect 7932 4496 7984 4505
rect 9128 4496 9180 4548
rect 9220 4496 9272 4548
rect 10324 4496 10376 4548
rect 6184 4428 6236 4480
rect 6552 4428 6604 4480
rect 10140 4428 10192 4480
rect 10508 4539 10560 4548
rect 10508 4505 10517 4539
rect 10517 4505 10551 4539
rect 10551 4505 10560 4539
rect 10508 4496 10560 4505
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 11060 4564 11112 4616
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 10692 4428 10744 4480
rect 2955 4326 3007 4378
rect 3019 4326 3071 4378
rect 3083 4326 3135 4378
rect 3147 4326 3199 4378
rect 3211 4326 3263 4378
rect 5646 4326 5698 4378
rect 5710 4326 5762 4378
rect 5774 4326 5826 4378
rect 5838 4326 5890 4378
rect 5902 4326 5954 4378
rect 8337 4326 8389 4378
rect 8401 4326 8453 4378
rect 8465 4326 8517 4378
rect 8529 4326 8581 4378
rect 8593 4326 8645 4378
rect 11028 4326 11080 4378
rect 11092 4326 11144 4378
rect 11156 4326 11208 4378
rect 11220 4326 11272 4378
rect 11284 4326 11336 4378
rect 3608 4224 3660 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2688 4156 2740 4208
rect 5540 4224 5592 4276
rect 7196 4224 7248 4276
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 7932 4224 7984 4276
rect 940 4020 992 4072
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 7104 4156 7156 4208
rect 2136 4020 2188 4072
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 2688 3884 2740 3936
rect 4712 4020 4764 4072
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6184 4088 6236 4140
rect 6276 4088 6328 4140
rect 8116 4131 8168 4140
rect 8116 4097 8161 4131
rect 8161 4097 8168 4131
rect 8116 4088 8168 4097
rect 8668 4088 8720 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 10784 4156 10836 4208
rect 9404 4088 9456 4097
rect 8024 4020 8076 4072
rect 10048 4020 10100 4072
rect 10324 4063 10376 4072
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 9036 3952 9088 4004
rect 9128 3952 9180 4004
rect 4804 3884 4856 3936
rect 5448 3884 5500 3936
rect 6276 3884 6328 3936
rect 6920 3884 6972 3936
rect 8116 3884 8168 3936
rect 11428 3952 11480 4004
rect 10232 3884 10284 3936
rect 2295 3782 2347 3834
rect 2359 3782 2411 3834
rect 2423 3782 2475 3834
rect 2487 3782 2539 3834
rect 2551 3782 2603 3834
rect 4986 3782 5038 3834
rect 5050 3782 5102 3834
rect 5114 3782 5166 3834
rect 5178 3782 5230 3834
rect 5242 3782 5294 3834
rect 7677 3782 7729 3834
rect 7741 3782 7793 3834
rect 7805 3782 7857 3834
rect 7869 3782 7921 3834
rect 7933 3782 7985 3834
rect 10368 3782 10420 3834
rect 10432 3782 10484 3834
rect 10496 3782 10548 3834
rect 10560 3782 10612 3834
rect 10624 3782 10676 3834
rect 2780 3680 2832 3732
rect 5448 3680 5500 3732
rect 6552 3680 6604 3732
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3608 3587 3660 3596
rect 3608 3553 3617 3587
rect 3617 3553 3651 3587
rect 3651 3553 3660 3587
rect 3608 3544 3660 3553
rect 5448 3544 5500 3596
rect 4252 3476 4304 3528
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 10232 3723 10284 3732
rect 10232 3689 10241 3723
rect 10241 3689 10275 3723
rect 10275 3689 10284 3723
rect 10232 3680 10284 3689
rect 7564 3612 7616 3664
rect 6184 3476 6236 3528
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 4804 3408 4856 3460
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7380 3451 7432 3460
rect 7380 3417 7389 3451
rect 7389 3417 7423 3451
rect 7423 3417 7432 3451
rect 7380 3408 7432 3417
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 6920 3340 6972 3392
rect 7472 3340 7524 3392
rect 8208 3408 8260 3460
rect 8760 3612 8812 3664
rect 8944 3544 8996 3596
rect 10692 3544 10744 3596
rect 8116 3340 8168 3392
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 2955 3238 3007 3290
rect 3019 3238 3071 3290
rect 3083 3238 3135 3290
rect 3147 3238 3199 3290
rect 3211 3238 3263 3290
rect 5646 3238 5698 3290
rect 5710 3238 5762 3290
rect 5774 3238 5826 3290
rect 5838 3238 5890 3290
rect 5902 3238 5954 3290
rect 8337 3238 8389 3290
rect 8401 3238 8453 3290
rect 8465 3238 8517 3290
rect 8529 3238 8581 3290
rect 8593 3238 8645 3290
rect 11028 3238 11080 3290
rect 11092 3238 11144 3290
rect 11156 3238 11208 3290
rect 11220 3238 11272 3290
rect 11284 3238 11336 3290
rect 2596 3136 2648 3188
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 4804 3136 4856 3188
rect 5356 3136 5408 3188
rect 6092 3136 6144 3188
rect 1676 3068 1728 3120
rect 7196 3136 7248 3188
rect 7472 3136 7524 3188
rect 1308 3000 1360 3052
rect 20 2932 72 2984
rect 3792 2932 3844 2984
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 5172 2932 5224 2984
rect 2320 2907 2372 2916
rect 2320 2873 2329 2907
rect 2329 2873 2363 2907
rect 2363 2873 2372 2907
rect 2320 2864 2372 2873
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5816 3000 5868 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 6460 3000 6512 3052
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7656 3000 7708 3052
rect 6184 2864 6236 2916
rect 6460 2907 6512 2916
rect 6460 2873 6469 2907
rect 6469 2873 6503 2907
rect 6503 2873 6512 2907
rect 6460 2864 6512 2873
rect 7656 2864 7708 2916
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 10048 3136 10100 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11612 3136 11664 3188
rect 10416 3068 10468 3120
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 8760 3043 8812 3052
rect 8760 3009 8768 3043
rect 8768 3009 8802 3043
rect 8802 3009 8812 3043
rect 8760 3000 8812 3009
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 11336 3043 11388 3052
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 8116 2864 8168 2916
rect 1492 2796 1544 2848
rect 6644 2796 6696 2848
rect 7380 2796 7432 2848
rect 7932 2796 7984 2848
rect 9036 2864 9088 2916
rect 2295 2694 2347 2746
rect 2359 2694 2411 2746
rect 2423 2694 2475 2746
rect 2487 2694 2539 2746
rect 2551 2694 2603 2746
rect 4986 2694 5038 2746
rect 5050 2694 5102 2746
rect 5114 2694 5166 2746
rect 5178 2694 5230 2746
rect 5242 2694 5294 2746
rect 7677 2694 7729 2746
rect 7741 2694 7793 2746
rect 7805 2694 7857 2746
rect 7869 2694 7921 2746
rect 7933 2694 7985 2746
rect 10368 2694 10420 2746
rect 10432 2694 10484 2746
rect 10496 2694 10548 2746
rect 10560 2694 10612 2746
rect 10624 2694 10676 2746
rect 5540 2592 5592 2644
rect 6460 2592 6512 2644
rect 7472 2592 7524 2644
rect 9956 2592 10008 2644
rect 10784 2592 10836 2644
rect 11428 2592 11480 2644
rect 7196 2524 7248 2576
rect 11520 2524 11572 2576
rect 1952 2456 2004 2508
rect 3608 2456 3660 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 7288 2456 7340 2508
rect 4896 2388 4948 2440
rect 5172 2388 5224 2440
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7196 2388 7248 2440
rect 7748 2388 7800 2440
rect 8116 2388 8168 2440
rect 11428 2456 11480 2508
rect 10416 2388 10468 2440
rect 3424 2320 3476 2372
rect 6460 2320 6512 2372
rect 11612 2388 11664 2440
rect 12900 2320 12952 2372
rect 4712 2252 4764 2304
rect 9036 2252 9088 2304
rect 2955 2150 3007 2202
rect 3019 2150 3071 2202
rect 3083 2150 3135 2202
rect 3147 2150 3199 2202
rect 3211 2150 3263 2202
rect 5646 2150 5698 2202
rect 5710 2150 5762 2202
rect 5774 2150 5826 2202
rect 5838 2150 5890 2202
rect 5902 2150 5954 2202
rect 8337 2150 8389 2202
rect 8401 2150 8453 2202
rect 8465 2150 8517 2202
rect 8529 2150 8581 2202
rect 8593 2150 8645 2202
rect 11028 2150 11080 2202
rect 11092 2150 11144 2202
rect 11156 2150 11208 2202
rect 11220 2150 11272 2202
rect 11284 2150 11336 2202
<< metal2 >>
rect 18 14397 74 15197
rect 1306 14397 1362 15197
rect 2594 14397 2650 15197
rect 3882 14397 3938 15197
rect 5170 14397 5226 15197
rect 6458 14498 6514 15197
rect 6458 14470 6592 14498
rect 6458 14397 6514 14470
rect 32 12306 60 14397
rect 1030 12336 1086 12345
rect 20 12300 72 12306
rect 1030 12271 1086 12280
rect 20 12242 72 12248
rect 1044 12238 1072 12271
rect 1032 12232 1084 12238
rect 1032 12174 1084 12180
rect 1320 11762 1348 14397
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1504 12442 1532 13631
rect 2608 13410 2636 14397
rect 2608 13382 2728 13410
rect 2295 12540 2603 12549
rect 2295 12538 2301 12540
rect 2357 12538 2381 12540
rect 2437 12538 2461 12540
rect 2517 12538 2541 12540
rect 2597 12538 2603 12540
rect 2357 12486 2359 12538
rect 2539 12486 2541 12538
rect 2295 12484 2301 12486
rect 2357 12484 2381 12486
rect 2437 12484 2461 12486
rect 2517 12484 2541 12486
rect 2597 12484 2603 12486
rect 2295 12475 2603 12484
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 2700 12238 2728 13382
rect 3896 12442 3924 14397
rect 5184 13274 5212 14397
rect 5184 13246 5396 13274
rect 4986 12540 5294 12549
rect 4986 12538 4992 12540
rect 5048 12538 5072 12540
rect 5128 12538 5152 12540
rect 5208 12538 5232 12540
rect 5288 12538 5294 12540
rect 5048 12486 5050 12538
rect 5230 12486 5232 12538
rect 4986 12484 4992 12486
rect 5048 12484 5072 12486
rect 5128 12484 5152 12486
rect 5208 12484 5232 12486
rect 5288 12484 5294 12486
rect 4986 12475 5294 12484
rect 5368 12442 5396 13246
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1780 11898 1808 12106
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 952 10674 980 10911
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1596 9382 1624 11494
rect 1688 11354 1716 11562
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1688 9654 1716 11290
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1688 8634 1716 9590
rect 1780 9586 1808 11834
rect 1860 11688 1912 11694
rect 1858 11656 1860 11665
rect 2688 11688 2740 11694
rect 1912 11656 1914 11665
rect 2688 11630 2740 11636
rect 1858 11591 1914 11600
rect 1872 11150 1900 11591
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 11286 1992 11494
rect 2295 11452 2603 11461
rect 2295 11450 2301 11452
rect 2357 11450 2381 11452
rect 2437 11450 2461 11452
rect 2517 11450 2541 11452
rect 2597 11450 2603 11452
rect 2357 11398 2359 11450
rect 2539 11398 2541 11450
rect 2295 11396 2301 11398
rect 2357 11396 2381 11398
rect 2437 11396 2461 11398
rect 2517 11396 2541 11398
rect 2597 11396 2603 11398
rect 2295 11387 2603 11396
rect 2700 11354 2728 11630
rect 2884 11558 2912 12038
rect 2955 11996 3263 12005
rect 2955 11994 2961 11996
rect 3017 11994 3041 11996
rect 3097 11994 3121 11996
rect 3177 11994 3201 11996
rect 3257 11994 3263 11996
rect 3017 11942 3019 11994
rect 3199 11942 3201 11994
rect 2955 11940 2961 11942
rect 3017 11940 3041 11942
rect 3097 11940 3121 11942
rect 3177 11940 3201 11942
rect 3257 11940 3263 11942
rect 2955 11931 3263 11940
rect 4080 11762 4108 12242
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4264 11830 4292 12174
rect 4528 11892 4580 11898
rect 4448 11852 4528 11880
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 10674 1992 10950
rect 2056 10810 2084 11290
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2240 10674 2268 11222
rect 2792 10742 2820 11222
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10810 2912 11086
rect 3436 11082 3464 11562
rect 3528 11286 3556 11562
rect 3884 11552 3936 11558
rect 3936 11500 4016 11506
rect 3884 11494 4016 11500
rect 3896 11478 4016 11494
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3528 11150 3556 11222
rect 3620 11150 3648 11290
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2955 10908 3263 10917
rect 2955 10906 2961 10908
rect 3017 10906 3041 10908
rect 3097 10906 3121 10908
rect 3177 10906 3201 10908
rect 3257 10906 3263 10908
rect 3017 10854 3019 10906
rect 3199 10854 3201 10906
rect 2955 10852 2961 10854
rect 3017 10852 3041 10854
rect 3097 10852 3121 10854
rect 3177 10852 3201 10854
rect 3257 10852 3263 10854
rect 2955 10843 3263 10852
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1872 10062 1900 10406
rect 2056 10062 2084 10406
rect 2295 10364 2603 10373
rect 2295 10362 2301 10364
rect 2357 10362 2381 10364
rect 2437 10362 2461 10364
rect 2517 10362 2541 10364
rect 2597 10362 2603 10364
rect 2357 10310 2359 10362
rect 2539 10310 2541 10362
rect 2295 10308 2301 10310
rect 2357 10308 2381 10310
rect 2437 10308 2461 10310
rect 2517 10308 2541 10310
rect 2597 10308 2603 10310
rect 2295 10299 2603 10308
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 8838 1808 9522
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1492 8288 1544 8294
rect 1398 8256 1454 8265
rect 1492 8230 1544 8236
rect 1398 8191 1454 8200
rect 1504 7886 1532 8230
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 1398 6896 1454 6905
rect 1504 6866 1532 7822
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6934 1624 7142
rect 1584 6928 1636 6934
rect 1584 6870 1636 6876
rect 1398 6831 1454 6840
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 5302 980 5471
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 1308 4480 1360 4486
rect 1308 4422 1360 4428
rect 1320 4185 1348 4422
rect 1306 4176 1362 4185
rect 1306 4111 1362 4120
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 20 2984 72 2990
rect 20 2926 72 2932
rect 32 800 60 2926
rect 952 2825 980 4014
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1320 800 1348 2994
rect 1412 1465 1440 4082
rect 1504 2854 1532 6802
rect 1688 5273 1716 8026
rect 1780 5778 1808 8774
rect 2056 8566 2084 9998
rect 2884 9586 2912 10474
rect 3344 10146 3372 10950
rect 3252 10118 3372 10146
rect 3436 10130 3464 11018
rect 3424 10124 3476 10130
rect 3252 10062 3280 10118
rect 3424 10066 3476 10072
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 2955 9820 3263 9829
rect 2955 9818 2961 9820
rect 3017 9818 3041 9820
rect 3097 9818 3121 9820
rect 3177 9818 3201 9820
rect 3257 9818 3263 9820
rect 3017 9766 3019 9818
rect 3199 9766 3201 9818
rect 2955 9764 2961 9766
rect 3017 9764 3041 9766
rect 3097 9764 3121 9766
rect 3177 9764 3201 9766
rect 3257 9764 3263 9766
rect 2955 9755 3263 9764
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2148 9042 2176 9318
rect 2295 9276 2603 9285
rect 2295 9274 2301 9276
rect 2357 9274 2381 9276
rect 2437 9274 2461 9276
rect 2517 9274 2541 9276
rect 2597 9274 2603 9276
rect 2357 9222 2359 9274
rect 2539 9222 2541 9274
rect 2295 9220 2301 9222
rect 2357 9220 2381 9222
rect 2437 9220 2461 9222
rect 2517 9220 2541 9222
rect 2597 9220 2603 9222
rect 2295 9211 2603 9220
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2148 8634 2176 8978
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2516 8566 2544 8910
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1674 5264 1730 5273
rect 1674 5199 1730 5208
rect 1582 4040 1638 4049
rect 1582 3975 1584 3984
rect 1636 3975 1638 3984
rect 1584 3946 1636 3952
rect 1688 3126 1716 5199
rect 1872 4010 1900 7278
rect 1964 5302 1992 7958
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7546 2084 7822
rect 2148 7750 2176 8434
rect 2295 8188 2603 8197
rect 2295 8186 2301 8188
rect 2357 8186 2381 8188
rect 2437 8186 2461 8188
rect 2517 8186 2541 8188
rect 2597 8186 2603 8188
rect 2357 8134 2359 8186
rect 2539 8134 2541 8186
rect 2295 8132 2301 8134
rect 2357 8132 2381 8134
rect 2437 8132 2461 8134
rect 2517 8132 2541 8134
rect 2597 8132 2603 8134
rect 2295 8123 2603 8132
rect 2596 8084 2648 8090
rect 2700 8072 2728 8978
rect 3252 8956 3280 9318
rect 3344 9110 3372 9998
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3528 9382 3556 9930
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3252 8928 3372 8956
rect 2955 8732 3263 8741
rect 2955 8730 2961 8732
rect 3017 8730 3041 8732
rect 3097 8730 3121 8732
rect 3177 8730 3201 8732
rect 3257 8730 3263 8732
rect 3017 8678 3019 8730
rect 3199 8678 3201 8730
rect 2955 8676 2961 8678
rect 3017 8676 3041 8678
rect 3097 8676 3121 8678
rect 3177 8676 3201 8678
rect 3257 8676 3263 8678
rect 2955 8667 3263 8676
rect 3344 8616 3372 8928
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3252 8588 3372 8616
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2648 8044 2728 8072
rect 2596 8026 2648 8032
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2240 7342 2268 7822
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7478 2360 7754
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2700 7410 2728 7686
rect 2792 7546 2820 8434
rect 3252 8022 3280 8588
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8016 3292 8022
rect 3238 7984 3240 7993
rect 3292 7984 3294 7993
rect 3238 7919 3294 7928
rect 3344 7868 3372 8434
rect 3436 7886 3464 8774
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 7954 3556 8366
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 2884 7840 3372 7868
rect 3424 7880 3476 7886
rect 2884 7750 2912 7840
rect 3424 7822 3476 7828
rect 3514 7848 3570 7857
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2955 7644 3263 7653
rect 2955 7642 2961 7644
rect 3017 7642 3041 7644
rect 3097 7642 3121 7644
rect 3177 7642 3201 7644
rect 3257 7642 3263 7644
rect 3017 7590 3019 7642
rect 3199 7590 3201 7642
rect 2955 7588 2961 7590
rect 3017 7588 3041 7590
rect 3097 7588 3121 7590
rect 3177 7588 3201 7590
rect 3257 7588 3263 7590
rect 2955 7579 3263 7588
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2976 7410 3004 7482
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 3436 7342 3464 7822
rect 3514 7783 3570 7792
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2295 7100 2603 7109
rect 2295 7098 2301 7100
rect 2357 7098 2381 7100
rect 2437 7098 2461 7100
rect 2517 7098 2541 7100
rect 2597 7098 2603 7100
rect 2357 7046 2359 7098
rect 2539 7046 2541 7098
rect 2295 7044 2301 7046
rect 2357 7044 2381 7046
rect 2437 7044 2461 7046
rect 2517 7044 2541 7046
rect 2597 7044 2603 7046
rect 2295 7035 2603 7044
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1964 2514 1992 5238
rect 2148 4078 2176 6258
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2295 6012 2603 6021
rect 2295 6010 2301 6012
rect 2357 6010 2381 6012
rect 2437 6010 2461 6012
rect 2517 6010 2541 6012
rect 2597 6010 2603 6012
rect 2357 5958 2359 6010
rect 2539 5958 2541 6010
rect 2295 5956 2301 5958
rect 2357 5956 2381 5958
rect 2437 5956 2461 5958
rect 2517 5956 2541 5958
rect 2597 5956 2603 5958
rect 2295 5947 2603 5956
rect 2700 5778 2728 6190
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5302 2728 5714
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2295 4924 2603 4933
rect 2295 4922 2301 4924
rect 2357 4922 2381 4924
rect 2437 4922 2461 4924
rect 2517 4922 2541 4924
rect 2597 4922 2603 4924
rect 2357 4870 2359 4922
rect 2539 4870 2541 4922
rect 2295 4868 2301 4870
rect 2357 4868 2381 4870
rect 2437 4868 2461 4870
rect 2517 4868 2541 4870
rect 2597 4868 2603 4870
rect 2295 4859 2603 4868
rect 2700 4706 2728 5238
rect 2608 4690 2728 4706
rect 2596 4684 2728 4690
rect 2648 4678 2728 4684
rect 2596 4626 2648 4632
rect 2700 4214 2728 4678
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2295 3836 2603 3845
rect 2295 3834 2301 3836
rect 2357 3834 2381 3836
rect 2437 3834 2461 3836
rect 2517 3834 2541 3836
rect 2597 3834 2603 3836
rect 2357 3782 2359 3834
rect 2539 3782 2541 3834
rect 2295 3780 2301 3782
rect 2357 3780 2381 3782
rect 2437 3780 2461 3782
rect 2517 3780 2541 3782
rect 2597 3780 2603 3782
rect 2295 3771 2603 3780
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2608 3097 2636 3130
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2318 2952 2374 2961
rect 2318 2887 2320 2896
rect 2372 2887 2374 2896
rect 2320 2858 2372 2864
rect 2295 2748 2603 2757
rect 2295 2746 2301 2748
rect 2357 2746 2381 2748
rect 2437 2746 2461 2748
rect 2517 2746 2541 2748
rect 2597 2746 2603 2748
rect 2357 2694 2359 2746
rect 2539 2694 2541 2746
rect 2295 2692 2301 2694
rect 2357 2692 2381 2694
rect 2437 2692 2461 2694
rect 2517 2692 2541 2694
rect 2597 2692 2603 2694
rect 2295 2683 2603 2692
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2700 2122 2728 3878
rect 2792 3738 2820 7142
rect 2955 6556 3263 6565
rect 2955 6554 2961 6556
rect 3017 6554 3041 6556
rect 3097 6554 3121 6556
rect 3177 6554 3201 6556
rect 3257 6554 3263 6556
rect 3017 6502 3019 6554
rect 3199 6502 3201 6554
rect 2955 6500 2961 6502
rect 3017 6500 3041 6502
rect 3097 6500 3121 6502
rect 3177 6500 3201 6502
rect 3257 6500 3263 6502
rect 2955 6491 3263 6500
rect 3528 6186 3556 7783
rect 3620 6225 3648 11086
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3804 10810 3832 11018
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 9110 3832 9454
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3804 7886 3832 9046
rect 3896 8566 3924 9590
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3712 7410 3740 7686
rect 3804 7478 3832 7822
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3804 6798 3832 7414
rect 3896 7206 3924 8026
rect 3988 7410 4016 11478
rect 4080 11082 4108 11698
rect 4448 11558 4476 11852
rect 4528 11834 4580 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4264 11121 4292 11494
rect 4250 11112 4306 11121
rect 4068 11076 4120 11082
rect 4250 11047 4252 11056
rect 4068 11018 4120 11024
rect 4304 11047 4306 11056
rect 4252 11018 4304 11024
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4172 10062 4200 10746
rect 4448 10146 4476 10950
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4356 10118 4476 10146
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9654 4200 9998
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4264 9586 4292 10066
rect 4356 10062 4384 10118
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 8974 4108 9318
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8090 4108 8910
rect 4172 8430 4200 9454
rect 4264 8498 4292 9522
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4080 7274 4108 7822
rect 4172 7750 4200 8366
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4264 7546 4292 7754
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 7478 4384 9998
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4448 9586 4476 9930
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4540 9466 4568 11698
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9586 4660 9862
rect 4724 9654 4752 11086
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10266 4844 11018
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4448 9438 4568 9466
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4448 7290 4476 9438
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4264 7262 4476 7290
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3896 7002 3924 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3988 6866 4016 7142
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3606 6216 3662 6225
rect 3516 6180 3568 6186
rect 3606 6151 3662 6160
rect 3516 6122 3568 6128
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 2955 5468 3263 5477
rect 2955 5466 2961 5468
rect 3017 5466 3041 5468
rect 3097 5466 3121 5468
rect 3177 5466 3201 5468
rect 3257 5466 3263 5468
rect 3017 5414 3019 5466
rect 3199 5414 3201 5466
rect 2955 5412 2961 5414
rect 3017 5412 3041 5414
rect 3097 5412 3121 5414
rect 3177 5412 3201 5414
rect 3257 5412 3263 5414
rect 2955 5403 3263 5412
rect 3330 4584 3386 4593
rect 3330 4519 3386 4528
rect 2955 4380 3263 4389
rect 2955 4378 2961 4380
rect 3017 4378 3041 4380
rect 3097 4378 3121 4380
rect 3177 4378 3201 4380
rect 3257 4378 3263 4380
rect 3017 4326 3019 4378
rect 3199 4326 3201 4378
rect 2955 4324 2961 4326
rect 3017 4324 3041 4326
rect 3097 4324 3121 4326
rect 3177 4324 3201 4326
rect 3257 4324 3263 4326
rect 2955 4315 3263 4324
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3344 3602 3372 4519
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 2955 3292 3263 3301
rect 2955 3290 2961 3292
rect 3017 3290 3041 3292
rect 3097 3290 3121 3292
rect 3177 3290 3201 3292
rect 3257 3290 3263 3292
rect 3017 3238 3019 3290
rect 3199 3238 3201 3290
rect 2955 3236 2961 3238
rect 3017 3236 3041 3238
rect 3097 3236 3121 3238
rect 3177 3236 3201 3238
rect 3257 3236 3263 3238
rect 2955 3227 3263 3236
rect 3436 2378 3464 6054
rect 4172 5710 4200 6598
rect 4264 5846 4292 7262
rect 4436 6928 4488 6934
rect 4540 6882 4568 9318
rect 4632 8906 4660 9522
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4816 8838 4844 9454
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8090 4660 8434
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4724 8022 4752 8502
rect 4712 8016 4764 8022
rect 4618 7984 4674 7993
rect 4712 7958 4764 7964
rect 4618 7919 4674 7928
rect 4488 6876 4568 6882
rect 4436 6870 4568 6876
rect 4448 6854 4568 6870
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4356 6458 4384 6666
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4540 6322 4568 6854
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3620 4282 3648 4490
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3620 2514 3648 3538
rect 4172 2990 4200 4966
rect 4356 4826 4384 6258
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4448 4146 4476 5782
rect 4632 5302 4660 7919
rect 4724 6254 4752 7958
rect 4816 7886 4844 8774
rect 4908 8294 4936 12310
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 4986 11452 5294 11461
rect 4986 11450 4992 11452
rect 5048 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5294 11452
rect 5048 11398 5050 11450
rect 5230 11398 5232 11450
rect 4986 11396 4992 11398
rect 5048 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5294 11398
rect 4986 11387 5294 11396
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5000 10742 5028 11222
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4986 10364 5294 10373
rect 4986 10362 4992 10364
rect 5048 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5294 10364
rect 5048 10310 5050 10362
rect 5230 10310 5232 10362
rect 4986 10308 4992 10310
rect 5048 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5294 10310
rect 4986 10299 5294 10308
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9382 5304 9930
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4986 9276 5294 9285
rect 4986 9274 4992 9276
rect 5048 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5294 9276
rect 5048 9222 5050 9274
rect 5230 9222 5232 9274
rect 4986 9220 4992 9222
rect 5048 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5294 9222
rect 4986 9211 5294 9220
rect 5368 8922 5396 12174
rect 5552 11830 5580 12378
rect 6564 12238 6592 14470
rect 7746 14397 7802 15197
rect 9034 14397 9090 15197
rect 10322 14397 10378 15197
rect 11610 14397 11666 15197
rect 12898 14397 12954 15197
rect 7760 12646 7788 14397
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 7677 12540 7985 12549
rect 7677 12538 7683 12540
rect 7739 12538 7763 12540
rect 7819 12538 7843 12540
rect 7899 12538 7923 12540
rect 7979 12538 7985 12540
rect 7739 12486 7741 12538
rect 7921 12486 7923 12538
rect 7677 12484 7683 12486
rect 7739 12484 7763 12486
rect 7819 12484 7843 12486
rect 7899 12484 7923 12486
rect 7979 12484 7985 12486
rect 7677 12475 7985 12484
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 5646 11996 5954 12005
rect 5646 11994 5652 11996
rect 5708 11994 5732 11996
rect 5788 11994 5812 11996
rect 5868 11994 5892 11996
rect 5948 11994 5954 11996
rect 5708 11942 5710 11994
rect 5890 11942 5892 11994
rect 5646 11940 5652 11942
rect 5708 11940 5732 11942
rect 5788 11940 5812 11942
rect 5868 11940 5892 11942
rect 5948 11940 5954 11942
rect 5646 11931 5954 11940
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5552 11336 5580 11766
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5460 11308 5580 11336
rect 5460 10062 5488 11308
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 11082 5580 11154
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10266 5580 11018
rect 5646 10908 5954 10917
rect 5646 10906 5652 10908
rect 5708 10906 5732 10908
rect 5788 10906 5812 10908
rect 5868 10906 5892 10908
rect 5948 10906 5954 10908
rect 5708 10854 5710 10906
rect 5890 10854 5892 10906
rect 5646 10852 5652 10854
rect 5708 10852 5732 10854
rect 5788 10852 5812 10854
rect 5868 10852 5892 10854
rect 5948 10852 5954 10854
rect 5646 10843 5954 10852
rect 6012 10606 6040 11630
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 10674 6132 11018
rect 6196 11014 6224 11562
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6104 10554 6132 10610
rect 6104 10538 6224 10554
rect 6104 10532 6236 10538
rect 6104 10526 6184 10532
rect 6184 10474 6236 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 6012 10062 6040 10406
rect 5448 10056 5500 10062
rect 6000 10056 6052 10062
rect 5500 10004 5580 10010
rect 5448 9998 5580 10004
rect 6000 9998 6052 10004
rect 5460 9982 5580 9998
rect 5552 9654 5580 9982
rect 5646 9820 5954 9829
rect 5646 9818 5652 9820
rect 5708 9818 5732 9820
rect 5788 9818 5812 9820
rect 5868 9818 5892 9820
rect 5948 9818 5954 9820
rect 5708 9766 5710 9818
rect 5890 9766 5892 9818
rect 5646 9764 5652 9766
rect 5708 9764 5732 9766
rect 5788 9764 5812 9766
rect 5868 9764 5892 9766
rect 5948 9764 5954 9766
rect 5646 9755 5954 9764
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5736 9382 5764 9522
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5184 8894 5396 8922
rect 5184 8401 5212 8894
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5276 8498 5304 8774
rect 5368 8498 5396 8774
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5170 8392 5226 8401
rect 5170 8327 5226 8336
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4908 7818 4936 8230
rect 4986 8188 5294 8197
rect 4986 8186 4992 8188
rect 5048 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5294 8188
rect 5048 8134 5050 8186
rect 5230 8134 5232 8186
rect 4986 8132 4992 8134
rect 5048 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5294 8134
rect 4986 8123 5294 8132
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 5000 7546 5028 7822
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4252 3528 4304 3534
rect 4250 3496 4252 3505
rect 4304 3496 4306 3505
rect 4250 3431 4306 3440
rect 4632 3194 4660 4558
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 2955 2204 3263 2213
rect 2955 2202 2961 2204
rect 3017 2202 3041 2204
rect 3097 2202 3121 2204
rect 3177 2202 3201 2204
rect 3257 2202 3263 2204
rect 3017 2150 3019 2202
rect 3199 2150 3201 2202
rect 2955 2148 2961 2150
rect 3017 2148 3041 2150
rect 3097 2148 3121 2150
rect 3177 2148 3201 2150
rect 3257 2148 3263 2150
rect 2955 2139 3263 2148
rect 2608 2094 2728 2122
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 2608 800 2636 2094
rect 3804 1578 3832 2926
rect 4724 2310 4752 4014
rect 4816 3942 4844 7414
rect 5000 7290 5028 7482
rect 4908 7262 5028 7290
rect 4908 6798 4936 7262
rect 4986 7100 5294 7109
rect 4986 7098 4992 7100
rect 5048 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5294 7100
rect 5048 7046 5050 7098
rect 5230 7046 5232 7098
rect 4986 7044 4992 7046
rect 5048 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5294 7046
rect 4986 7035 5294 7044
rect 5368 6934 5396 7958
rect 5460 7886 5488 9114
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7206 5488 7822
rect 5552 7290 5580 9318
rect 6196 8974 6224 9522
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6196 8838 6224 8910
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6288 8786 6316 12106
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6472 11665 6500 11766
rect 6458 11656 6514 11665
rect 6458 11591 6514 11600
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11150 6408 11494
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6472 9602 6500 11591
rect 6380 9574 6500 9602
rect 6564 9586 6592 12038
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 9580 6604 9586
rect 6380 8945 6408 9574
rect 6552 9522 6604 9528
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6366 8936 6422 8945
rect 6366 8871 6422 8880
rect 5646 8732 5954 8741
rect 5646 8730 5652 8732
rect 5708 8730 5732 8732
rect 5788 8730 5812 8732
rect 5868 8730 5892 8732
rect 5948 8730 5954 8732
rect 5708 8678 5710 8730
rect 5890 8678 5892 8730
rect 5646 8676 5652 8678
rect 5708 8676 5732 8678
rect 5788 8676 5812 8678
rect 5868 8676 5892 8678
rect 5948 8676 5954 8678
rect 5646 8667 5954 8676
rect 6196 8650 6224 8774
rect 6288 8758 6408 8786
rect 6000 8628 6052 8634
rect 6196 8622 6316 8650
rect 6000 8570 6052 8576
rect 6012 8498 6040 8570
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5920 8378 5948 8434
rect 5920 8350 6040 8378
rect 6012 7750 6040 8350
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6104 8090 6132 8298
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5646 7644 5954 7653
rect 5646 7642 5652 7644
rect 5708 7642 5732 7644
rect 5788 7642 5812 7644
rect 5868 7642 5892 7644
rect 5948 7642 5954 7644
rect 5708 7590 5710 7642
rect 5890 7590 5892 7642
rect 5646 7588 5652 7590
rect 5708 7588 5732 7590
rect 5788 7588 5812 7590
rect 5868 7588 5892 7590
rect 5948 7588 5954 7590
rect 5646 7579 5954 7588
rect 6012 7478 6040 7686
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6000 7336 6052 7342
rect 5552 7262 5672 7290
rect 6000 7278 6052 7284
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5460 7002 5488 7142
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5000 6458 5028 6734
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5276 6322 5304 6598
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4986 6012 5294 6021
rect 4986 6010 4992 6012
rect 5048 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5294 6012
rect 5048 5958 5050 6010
rect 5230 5958 5232 6010
rect 4986 5956 4992 5958
rect 5048 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5294 5958
rect 4986 5947 5294 5956
rect 5368 5914 5396 6258
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5460 5846 5488 6054
rect 5552 5846 5580 7142
rect 5644 6866 5672 7262
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 6012 6798 6040 7278
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5736 6644 5764 6734
rect 5736 6616 6040 6644
rect 5646 6556 5954 6565
rect 5646 6554 5652 6556
rect 5708 6554 5732 6556
rect 5788 6554 5812 6556
rect 5868 6554 5892 6556
rect 5948 6554 5954 6556
rect 5708 6502 5710 6554
rect 5890 6502 5892 6554
rect 5646 6500 5652 6502
rect 5708 6500 5732 6502
rect 5788 6500 5812 6502
rect 5868 6500 5892 6502
rect 5948 6500 5954 6502
rect 5646 6491 5954 6500
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5828 6322 5856 6394
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5644 6089 5672 6190
rect 5630 6080 5686 6089
rect 5630 6015 5686 6024
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5828 5710 5856 6258
rect 5920 6186 5948 6258
rect 6012 6186 6040 6616
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6104 5642 6132 6870
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5448 5296 5500 5302
rect 5446 5264 5448 5273
rect 5500 5264 5502 5273
rect 5552 5250 5580 5510
rect 5646 5468 5954 5477
rect 5646 5466 5652 5468
rect 5708 5466 5732 5468
rect 5788 5466 5812 5468
rect 5868 5466 5892 5468
rect 5948 5466 5954 5468
rect 5708 5414 5710 5466
rect 5890 5414 5892 5466
rect 5646 5412 5652 5414
rect 5708 5412 5732 5414
rect 5788 5412 5812 5414
rect 5868 5412 5892 5414
rect 5948 5412 5954 5414
rect 5646 5403 5954 5412
rect 5552 5222 5948 5250
rect 6012 5234 6040 5510
rect 5446 5199 5502 5208
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5368 4978 5396 5034
rect 5368 4950 5580 4978
rect 4986 4924 5294 4933
rect 4986 4922 4992 4924
rect 5048 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5294 4924
rect 5048 4870 5050 4922
rect 5230 4870 5232 4922
rect 4986 4868 4992 4870
rect 5048 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5294 4870
rect 4986 4859 5294 4868
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4816 3194 4844 3402
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 2446 4936 4762
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4986 3836 5294 3845
rect 4986 3834 4992 3836
rect 5048 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5294 3836
rect 5048 3782 5050 3834
rect 5230 3782 5232 3834
rect 4986 3780 4992 3782
rect 5048 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5294 3782
rect 4986 3771 5294 3780
rect 5368 3194 5396 4558
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5460 3942 5488 4490
rect 5552 4282 5580 4950
rect 5814 4720 5870 4729
rect 5920 4706 5948 5222
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5920 4678 6040 4706
rect 5814 4655 5870 4664
rect 5828 4604 5856 4655
rect 5908 4616 5960 4622
rect 5828 4576 5908 4604
rect 5908 4558 5960 4564
rect 5646 4380 5954 4389
rect 5646 4378 5652 4380
rect 5708 4378 5732 4380
rect 5788 4378 5812 4380
rect 5868 4378 5892 4380
rect 5948 4378 5954 4380
rect 5708 4326 5710 4378
rect 5890 4326 5892 4378
rect 5646 4324 5652 4326
rect 5708 4324 5732 4326
rect 5788 4324 5812 4326
rect 5868 4324 5892 4326
rect 5948 4324 5954 4326
rect 5646 4315 5954 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 6012 4146 6040 4678
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3738 5488 3878
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5172 2984 5224 2990
rect 5460 2938 5488 3538
rect 5646 3292 5954 3301
rect 5646 3290 5652 3292
rect 5708 3290 5732 3292
rect 5788 3290 5812 3292
rect 5868 3290 5892 3292
rect 5948 3290 5954 3292
rect 5708 3238 5710 3290
rect 5890 3238 5892 3290
rect 5646 3236 5652 3238
rect 5708 3236 5732 3238
rect 5788 3236 5812 3238
rect 5868 3236 5892 3238
rect 5948 3236 5954 3238
rect 5646 3227 5954 3236
rect 6104 3194 6132 5170
rect 6196 4758 6224 8502
rect 6288 5710 6316 8622
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6380 5273 6408 8758
rect 6472 8022 6500 9454
rect 6564 8838 6592 9522
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6656 8634 6684 10066
rect 6748 9178 6776 12038
rect 7300 11762 7328 12174
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7116 11150 7144 11562
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10538 7052 11018
rect 7116 10674 7144 11086
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6564 8294 6592 8434
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6656 7886 6684 8570
rect 6748 8498 6776 8774
rect 6840 8566 6868 9930
rect 6932 9586 6960 10406
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6734 8392 6790 8401
rect 6932 8378 6960 9522
rect 7024 9382 7052 9522
rect 7208 9518 7236 10950
rect 7392 10810 7420 11630
rect 7576 11558 7604 12310
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7852 11558 7880 12242
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11762 7972 12038
rect 8036 11762 8064 12242
rect 8680 12238 8708 12582
rect 9048 12238 9076 14397
rect 10336 12730 10364 14397
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 10244 12702 10364 12730
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8300 12096 8352 12102
rect 8220 12056 8300 12084
rect 8220 11762 8248 12056
rect 8300 12038 8352 12044
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 8337 11996 8645 12005
rect 8337 11994 8343 11996
rect 8399 11994 8423 11996
rect 8479 11994 8503 11996
rect 8559 11994 8583 11996
rect 8639 11994 8645 11996
rect 8399 11942 8401 11994
rect 8581 11942 8583 11994
rect 8337 11940 8343 11942
rect 8399 11940 8423 11942
rect 8479 11940 8503 11942
rect 8559 11940 8583 11942
rect 8639 11940 8645 11942
rect 8337 11931 8645 11940
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7484 11150 7512 11222
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7300 10062 7328 10202
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 9722 7328 9862
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 9382 7236 9454
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7300 8566 7328 9658
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6734 8327 6790 8336
rect 6840 8350 6960 8378
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6748 7834 6776 8327
rect 6840 7954 6868 8350
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7886 6960 8230
rect 7024 7886 7052 8434
rect 6920 7880 6972 7886
rect 6656 7410 6684 7822
rect 6748 7806 6868 7834
rect 6920 7822 6972 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6564 6866 6592 7346
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6366 5264 6422 5273
rect 6366 5199 6422 5208
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6380 4690 6408 5199
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6182 4584 6238 4593
rect 6182 4519 6238 4528
rect 6196 4486 6224 4519
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6196 3913 6224 4082
rect 6288 4049 6316 4082
rect 6274 4040 6330 4049
rect 6274 3975 6330 3984
rect 6276 3936 6328 3942
rect 6182 3904 6238 3913
rect 6276 3878 6328 3884
rect 6182 3839 6238 3848
rect 6196 3534 6224 3839
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5814 3088 5870 3097
rect 5540 3052 5592 3058
rect 5814 3023 5816 3032
rect 5540 2994 5592 3000
rect 5868 3023 5870 3032
rect 5816 2994 5868 3000
rect 5224 2932 5488 2938
rect 5172 2926 5488 2932
rect 5184 2910 5488 2926
rect 4986 2748 5294 2757
rect 4986 2746 4992 2748
rect 5048 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5294 2748
rect 5048 2694 5050 2746
rect 5230 2694 5232 2746
rect 4986 2692 4992 2694
rect 5048 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5294 2694
rect 4986 2683 5294 2692
rect 5460 2514 5488 2910
rect 5552 2650 5580 2994
rect 5906 2952 5962 2961
rect 6196 2922 6224 3470
rect 6288 3040 6316 3878
rect 6380 3176 6408 4626
rect 6472 3534 6500 6666
rect 6734 6080 6790 6089
rect 6734 6015 6790 6024
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6564 4622 6592 5102
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 3738 6592 4422
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 3369 6500 3470
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6380 3148 6500 3176
rect 6472 3058 6500 3148
rect 6368 3052 6420 3058
rect 6288 3012 6368 3040
rect 6368 2994 6420 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6380 2961 6408 2994
rect 6366 2952 6422 2961
rect 5906 2887 5962 2896
rect 6184 2916 6236 2922
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5920 2446 5948 2887
rect 6366 2887 6422 2896
rect 6460 2916 6512 2922
rect 6184 2858 6236 2864
rect 6460 2858 6512 2864
rect 6472 2650 6500 2858
rect 6656 2854 6684 5646
rect 6748 3641 6776 6015
rect 6840 5642 6868 7806
rect 7116 7750 7144 8502
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7954 7236 8230
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6734 3632 6790 3641
rect 6734 3567 6790 3576
rect 6748 3534 6776 3567
rect 6736 3528 6788 3534
rect 6840 3505 6868 5578
rect 6932 5386 6960 7686
rect 7392 7342 7420 10746
rect 7484 10538 7512 11086
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7576 10010 7604 11494
rect 7677 11452 7985 11461
rect 7677 11450 7683 11452
rect 7739 11450 7763 11452
rect 7819 11450 7843 11452
rect 7899 11450 7923 11452
rect 7979 11450 7985 11452
rect 7739 11398 7741 11450
rect 7921 11398 7923 11450
rect 7677 11396 7683 11398
rect 7739 11396 7763 11398
rect 7819 11396 7843 11398
rect 7899 11396 7923 11398
rect 7979 11396 7985 11398
rect 7677 11387 7985 11396
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7944 11150 7972 11290
rect 8772 11150 8800 11494
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8760 11144 8812 11150
rect 8956 11121 8984 11562
rect 8760 11086 8812 11092
rect 8942 11112 8998 11121
rect 7944 10810 7972 11086
rect 8337 10908 8645 10917
rect 8337 10906 8343 10908
rect 8399 10906 8423 10908
rect 8479 10906 8503 10908
rect 8559 10906 8583 10908
rect 8639 10906 8645 10908
rect 8399 10854 8401 10906
rect 8581 10854 8583 10906
rect 8337 10852 8343 10854
rect 8399 10852 8423 10854
rect 8479 10852 8503 10854
rect 8559 10852 8583 10854
rect 8639 10852 8645 10854
rect 8337 10843 8645 10852
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8772 10742 8800 11086
rect 8942 11047 8998 11056
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7677 10364 7985 10373
rect 7677 10362 7683 10364
rect 7739 10362 7763 10364
rect 7819 10362 7843 10364
rect 7899 10362 7923 10364
rect 7979 10362 7985 10364
rect 7739 10310 7741 10362
rect 7921 10310 7923 10362
rect 7677 10308 7683 10310
rect 7739 10308 7763 10310
rect 7819 10308 7843 10310
rect 7899 10308 7923 10310
rect 7979 10308 7985 10310
rect 7677 10299 7985 10308
rect 7484 9994 7604 10010
rect 7472 9988 7604 9994
rect 7524 9982 7604 9988
rect 7472 9930 7524 9936
rect 7484 9897 7512 9930
rect 7840 9920 7892 9926
rect 7470 9888 7526 9897
rect 7840 9862 7892 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7470 9823 7526 9832
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7484 9586 7512 9658
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7852 9450 7880 9862
rect 8036 9722 8064 9862
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7677 9276 7985 9285
rect 7677 9274 7683 9276
rect 7739 9274 7763 9276
rect 7819 9274 7843 9276
rect 7899 9274 7923 9276
rect 7979 9274 7985 9276
rect 7739 9222 7741 9274
rect 7921 9222 7923 9274
rect 7677 9220 7683 9222
rect 7739 9220 7763 9222
rect 7819 9220 7843 9222
rect 7899 9220 7923 9222
rect 7979 9220 7985 9222
rect 7677 9211 7985 9220
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7944 8634 7972 9046
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6390 7052 6598
rect 7484 6390 7512 7958
rect 7576 7546 7604 8230
rect 7677 8188 7985 8197
rect 7677 8186 7683 8188
rect 7739 8186 7763 8188
rect 7819 8186 7843 8188
rect 7899 8186 7923 8188
rect 7979 8186 7985 8188
rect 7739 8134 7741 8186
rect 7921 8134 7923 8186
rect 7677 8132 7683 8134
rect 7739 8132 7763 8134
rect 7819 8132 7843 8134
rect 7899 8132 7923 8134
rect 7979 8132 7985 8134
rect 7677 8123 7985 8132
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7677 7100 7985 7109
rect 7677 7098 7683 7100
rect 7739 7098 7763 7100
rect 7819 7098 7843 7100
rect 7899 7098 7923 7100
rect 7979 7098 7985 7100
rect 7739 7046 7741 7098
rect 7921 7046 7923 7098
rect 7677 7044 7683 7046
rect 7739 7044 7763 7046
rect 7819 7044 7843 7046
rect 7899 7044 7923 7046
rect 7979 7044 7985 7046
rect 7677 7035 7985 7044
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7012 6384 7064 6390
rect 7472 6384 7524 6390
rect 7012 6326 7064 6332
rect 7102 6352 7158 6361
rect 7024 5710 7052 6326
rect 7102 6287 7104 6296
rect 7156 6287 7158 6296
rect 7300 6332 7472 6338
rect 7300 6326 7524 6332
rect 7300 6310 7512 6326
rect 7668 6322 7696 6598
rect 7656 6316 7708 6322
rect 7104 6258 7156 6264
rect 7300 6118 7328 6310
rect 7656 6258 7708 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7654 6216 7710 6225
rect 7392 6118 7420 6190
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7380 6112 7432 6118
rect 7432 6072 7512 6100
rect 7380 6054 7432 6060
rect 7300 5778 7328 6054
rect 7288 5772 7340 5778
rect 7208 5732 7288 5760
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5574 7052 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6932 5358 7052 5386
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4729 6960 5238
rect 6918 4720 6974 4729
rect 6918 4655 6974 4664
rect 6932 4554 6960 4655
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6920 3936 6972 3942
rect 7024 3924 7052 5358
rect 7208 5302 7236 5732
rect 7288 5714 7340 5720
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7196 5296 7248 5302
rect 7300 5273 7328 5510
rect 7196 5238 7248 5244
rect 7286 5264 7342 5273
rect 7286 5199 7288 5208
rect 7340 5199 7342 5208
rect 7288 5170 7340 5176
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4758 7236 5034
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7208 4282 7236 4694
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6972 3896 7052 3924
rect 6920 3878 6972 3884
rect 6736 3470 6788 3476
rect 6826 3496 6882 3505
rect 6826 3431 6882 3440
rect 6932 3398 6960 3878
rect 7116 3754 7144 4150
rect 7024 3726 7144 3754
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 7024 2774 7052 3726
rect 7300 3720 7328 5170
rect 7392 4622 7420 5510
rect 7484 5166 7512 6072
rect 7576 5710 7604 6190
rect 7654 6151 7656 6160
rect 7708 6151 7710 6160
rect 7656 6122 7708 6128
rect 7677 6012 7985 6021
rect 7677 6010 7683 6012
rect 7739 6010 7763 6012
rect 7819 6010 7843 6012
rect 7899 6010 7923 6012
rect 7979 6010 7985 6012
rect 7739 5958 7741 6010
rect 7921 5958 7923 6010
rect 7677 5956 7683 5958
rect 7739 5956 7763 5958
rect 7819 5956 7843 5958
rect 7899 5956 7923 5958
rect 7979 5956 7985 5958
rect 7677 5947 7985 5956
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 5302 7604 5646
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7677 4924 7985 4933
rect 7677 4922 7683 4924
rect 7739 4922 7763 4924
rect 7819 4922 7843 4924
rect 7899 4922 7923 4924
rect 7979 4922 7985 4924
rect 7739 4870 7741 4922
rect 7921 4870 7923 4922
rect 7677 4868 7683 4870
rect 7739 4868 7763 4870
rect 7819 4868 7843 4870
rect 7899 4868 7923 4870
rect 7979 4868 7985 4870
rect 7677 4859 7985 4868
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7668 4282 7696 4762
rect 7932 4752 7984 4758
rect 7838 4720 7894 4729
rect 8036 4729 8064 9318
rect 8128 9110 8156 10406
rect 8220 10062 8248 10678
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10266 8340 10406
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8337 9820 8645 9829
rect 8337 9818 8343 9820
rect 8399 9818 8423 9820
rect 8479 9818 8503 9820
rect 8559 9818 8583 9820
rect 8639 9818 8645 9820
rect 8399 9766 8401 9818
rect 8581 9766 8583 9818
rect 8337 9764 8343 9766
rect 8399 9764 8423 9766
rect 8479 9764 8503 9766
rect 8559 9764 8583 9766
rect 8639 9764 8645 9766
rect 8337 9755 8645 9764
rect 8956 9586 8984 11047
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8220 8974 8248 9522
rect 8312 9178 8340 9522
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8680 8974 8708 9318
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7932 4694 7984 4700
rect 8022 4720 8078 4729
rect 7838 4655 7894 4664
rect 7852 4622 7880 4655
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7944 4554 7972 4694
rect 8022 4655 8078 4664
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7944 4282 7972 4490
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8128 4146 8156 8774
rect 8220 8514 8248 8910
rect 8337 8732 8645 8741
rect 8337 8730 8343 8732
rect 8399 8730 8423 8732
rect 8479 8730 8503 8732
rect 8559 8730 8583 8732
rect 8639 8730 8645 8732
rect 8399 8678 8401 8730
rect 8581 8678 8583 8730
rect 8337 8676 8343 8678
rect 8399 8676 8423 8678
rect 8479 8676 8503 8678
rect 8559 8676 8583 8678
rect 8639 8676 8645 8678
rect 8337 8667 8645 8676
rect 8772 8634 8800 9454
rect 8864 8974 8892 9522
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 9178 9076 9386
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8220 8486 8340 8514
rect 8312 7954 8340 8486
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8496 7886 8524 8570
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8772 7834 8800 8570
rect 8864 7954 8892 8910
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8956 8498 8984 8570
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8265 8984 8434
rect 8942 8256 8998 8265
rect 8942 8191 8998 8200
rect 9048 8022 9076 9114
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7834 8984 7890
rect 8772 7806 8984 7834
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8220 6458 8248 7686
rect 8337 7644 8645 7653
rect 8337 7642 8343 7644
rect 8399 7642 8423 7644
rect 8479 7642 8503 7644
rect 8559 7642 8583 7644
rect 8639 7642 8645 7644
rect 8399 7590 8401 7642
rect 8581 7590 8583 7642
rect 8337 7588 8343 7590
rect 8399 7588 8423 7590
rect 8479 7588 8503 7590
rect 8559 7588 8583 7590
rect 8639 7588 8645 7590
rect 8337 7579 8645 7588
rect 8337 6556 8645 6565
rect 8337 6554 8343 6556
rect 8399 6554 8423 6556
rect 8479 6554 8503 6556
rect 8559 6554 8583 6556
rect 8639 6554 8645 6556
rect 8399 6502 8401 6554
rect 8581 6502 8583 6554
rect 8337 6500 8343 6502
rect 8399 6500 8423 6502
rect 8479 6500 8503 6502
rect 8559 6500 8583 6502
rect 8639 6500 8645 6502
rect 8337 6491 8645 6500
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8298 6352 8354 6361
rect 8680 6322 8708 7686
rect 8772 6866 8800 7806
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8298 6287 8300 6296
rect 8352 6287 8354 6296
rect 8484 6316 8536 6322
rect 8300 6258 8352 6264
rect 8484 6258 8536 6264
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5302 8248 5714
rect 8312 5710 8340 6258
rect 8496 5778 8524 6258
rect 8956 5778 8984 6734
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8337 5468 8645 5477
rect 8337 5466 8343 5468
rect 8399 5466 8423 5468
rect 8479 5466 8503 5468
rect 8559 5466 8583 5468
rect 8639 5466 8645 5468
rect 8399 5414 8401 5466
rect 8581 5414 8583 5466
rect 8337 5412 8343 5414
rect 8399 5412 8423 5414
rect 8479 5412 8503 5414
rect 8559 5412 8583 5414
rect 8639 5412 8645 5414
rect 8337 5403 8645 5412
rect 8680 5352 8708 5646
rect 8496 5324 8708 5352
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8220 4758 8248 5238
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8496 4622 8524 5324
rect 8574 5264 8630 5273
rect 8630 5208 8892 5216
rect 8574 5199 8576 5208
rect 8628 5188 8892 5208
rect 8576 5170 8628 5176
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 4072 8076 4078
rect 8220 4026 8248 4558
rect 8337 4380 8645 4389
rect 8337 4378 8343 4380
rect 8399 4378 8423 4380
rect 8479 4378 8503 4380
rect 8559 4378 8583 4380
rect 8639 4378 8645 4380
rect 8399 4326 8401 4378
rect 8581 4326 8583 4378
rect 8337 4324 8343 4326
rect 8399 4324 8423 4326
rect 8479 4324 8503 4326
rect 8559 4324 8583 4326
rect 8639 4324 8645 4326
rect 8337 4315 8645 4324
rect 8680 4146 8708 4966
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8076 4020 8248 4026
rect 8024 4014 8248 4020
rect 8036 3998 8248 4014
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7677 3836 7985 3845
rect 7677 3834 7683 3836
rect 7739 3834 7763 3836
rect 7819 3834 7843 3836
rect 7899 3834 7923 3836
rect 7979 3834 7985 3836
rect 7739 3782 7741 3834
rect 7921 3782 7923 3834
rect 7677 3780 7683 3782
rect 7739 3780 7763 3782
rect 7819 3780 7843 3782
rect 7899 3780 7923 3782
rect 7979 3780 7985 3782
rect 7677 3771 7985 3780
rect 7208 3692 7328 3720
rect 7102 3632 7158 3641
rect 7102 3567 7158 3576
rect 7116 3534 7144 3567
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7208 3194 7236 3692
rect 7564 3664 7616 3670
rect 7300 3624 7564 3652
rect 7300 3534 7328 3624
rect 7564 3606 7616 3612
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6932 2746 7052 2774
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6932 2446 6960 2746
rect 7208 2582 7236 2994
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7208 2446 7236 2518
rect 7300 2514 7328 3470
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 3369 7420 3402
rect 7472 3392 7524 3398
rect 7378 3360 7434 3369
rect 7472 3334 7524 3340
rect 7378 3295 7434 3304
rect 7484 3194 7512 3334
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7484 3058 7512 3130
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7392 2854 7420 2994
rect 7668 2922 7696 2994
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7944 2854 7972 3470
rect 8128 3398 8156 3878
rect 8220 3602 8248 3998
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8220 3058 8248 3402
rect 8337 3292 8645 3301
rect 8337 3290 8343 3292
rect 8399 3290 8423 3292
rect 8479 3290 8503 3292
rect 8559 3290 8583 3292
rect 8639 3290 8645 3292
rect 8399 3238 8401 3290
rect 8581 3238 8583 3290
rect 8337 3236 8343 3238
rect 8399 3236 8423 3238
rect 8479 3236 8503 3238
rect 8559 3236 8583 3238
rect 8639 3236 8645 3238
rect 8337 3227 8645 3236
rect 8772 3058 8800 3606
rect 8864 3194 8892 5188
rect 8956 3602 8984 5714
rect 9048 4826 9076 7482
rect 9140 6390 9168 12038
rect 9416 11558 9444 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9232 8634 9260 9590
rect 9324 8838 9352 10134
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8906 9628 9318
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9324 8566 9352 8774
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8378 9444 8434
rect 9220 8356 9272 8362
rect 9416 8350 9536 8378
rect 9220 8298 9272 8304
rect 9232 8022 9260 8298
rect 9508 8294 9536 8350
rect 9312 8288 9364 8294
rect 9496 8288 9548 8294
rect 9312 8230 9364 8236
rect 9402 8256 9458 8265
rect 9324 8022 9352 8230
rect 9496 8230 9548 8236
rect 9402 8191 9458 8200
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9140 4672 9168 6326
rect 9232 6322 9260 7822
rect 9416 6798 9444 8191
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9324 6390 9352 6734
rect 9508 6730 9536 8230
rect 9600 8090 9628 8842
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9600 7750 9628 8026
rect 9692 7954 9720 11834
rect 9784 11150 9812 12310
rect 10244 12238 10272 12702
rect 10368 12540 10676 12549
rect 10368 12538 10374 12540
rect 10430 12538 10454 12540
rect 10510 12538 10534 12540
rect 10590 12538 10614 12540
rect 10670 12538 10676 12540
rect 10430 12486 10432 12538
rect 10612 12486 10614 12538
rect 10368 12484 10374 12486
rect 10430 12484 10454 12486
rect 10510 12484 10534 12486
rect 10590 12484 10614 12486
rect 10670 12484 10676 12486
rect 10368 12475 10676 12484
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9784 9110 9812 9522
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9784 8906 9812 9046
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9876 8294 9904 11698
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10470 9996 10542
rect 10060 10538 10088 12106
rect 10888 11762 10916 12106
rect 11028 11996 11336 12005
rect 11028 11994 11034 11996
rect 11090 11994 11114 11996
rect 11170 11994 11194 11996
rect 11250 11994 11274 11996
rect 11330 11994 11336 11996
rect 11090 11942 11092 11994
rect 11272 11942 11274 11994
rect 11028 11940 11034 11942
rect 11090 11940 11114 11942
rect 11170 11940 11194 11942
rect 11250 11940 11274 11942
rect 11330 11940 11336 11942
rect 11028 11931 11336 11940
rect 11440 11830 11468 13631
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11532 11694 11560 12271
rect 11624 11898 11652 14397
rect 12912 12442 12940 14397
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 10368 11452 10676 11461
rect 10368 11450 10374 11452
rect 10430 11450 10454 11452
rect 10510 11450 10534 11452
rect 10590 11450 10614 11452
rect 10670 11450 10676 11452
rect 10430 11398 10432 11450
rect 10612 11398 10614 11450
rect 10368 11396 10374 11398
rect 10430 11396 10454 11398
rect 10510 11396 10534 11398
rect 10590 11396 10614 11398
rect 10670 11396 10676 11398
rect 10368 11387 10676 11396
rect 10416 11348 10468 11354
rect 10244 11308 10416 11336
rect 10244 10742 10272 11308
rect 10416 11290 10468 11296
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10612 11150 10640 11222
rect 10888 11150 10916 11290
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9874 9996 10406
rect 10060 9994 10088 10474
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9968 9846 10088 9874
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 9110 9996 9318
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8498 9996 8910
rect 10060 8498 10088 9846
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7002 9628 7686
rect 9692 7002 9720 7890
rect 9876 7546 9904 8230
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6882 9812 7346
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9692 6854 9812 6882
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9232 5710 9260 6054
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9324 5302 9352 6054
rect 9508 5914 9536 6122
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5642 9628 6734
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9692 5030 9720 6854
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6322 9812 6598
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9140 4644 9260 4672
rect 9232 4554 9260 4644
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9140 4010 9168 4490
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8114 2952 8170 2961
rect 9048 2922 9076 3946
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 3641 9168 3674
rect 9126 3632 9182 3641
rect 9126 3567 9182 3576
rect 9416 3505 9444 4082
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9508 3058 9536 4762
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 3097 9720 4626
rect 9876 4049 9904 7142
rect 9862 4040 9918 4049
rect 9862 3975 9918 3984
rect 9678 3088 9734 3097
rect 9496 3052 9548 3058
rect 9678 3023 9734 3032
rect 9496 2994 9548 3000
rect 8114 2887 8116 2896
rect 8168 2887 8170 2896
rect 9036 2916 9088 2922
rect 8116 2858 8168 2864
rect 9036 2858 9088 2864
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7677 2748 7985 2757
rect 7677 2746 7683 2748
rect 7739 2746 7763 2748
rect 7819 2746 7843 2748
rect 7899 2746 7923 2748
rect 7979 2746 7985 2748
rect 7739 2694 7741 2746
rect 7921 2694 7923 2746
rect 7677 2692 7683 2694
rect 7739 2692 7763 2694
rect 7819 2692 7843 2694
rect 7899 2692 7923 2694
rect 7979 2692 7985 2694
rect 7470 2680 7526 2689
rect 7677 2683 7985 2692
rect 7470 2615 7472 2624
rect 7524 2615 7526 2624
rect 7472 2586 7524 2592
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 8128 2446 8156 2858
rect 9968 2650 9996 8434
rect 10060 6905 10088 8434
rect 10046 6896 10102 6905
rect 10046 6831 10102 6840
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6458 10088 6598
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 5914 10088 6394
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10152 5642 10180 10474
rect 10244 10198 10272 10678
rect 10612 10538 10640 11086
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10368 10364 10676 10373
rect 10368 10362 10374 10364
rect 10430 10362 10454 10364
rect 10510 10362 10534 10364
rect 10590 10362 10614 10364
rect 10670 10362 10676 10364
rect 10430 10310 10432 10362
rect 10612 10310 10614 10362
rect 10368 10308 10374 10310
rect 10430 10308 10454 10310
rect 10510 10308 10534 10310
rect 10590 10308 10614 10310
rect 10670 10308 10676 10310
rect 10368 10299 10676 10308
rect 10704 10266 10732 11018
rect 10796 10810 10824 11018
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 10674 10916 11086
rect 11532 10985 11560 11086
rect 11518 10976 11574 10985
rect 11028 10908 11336 10917
rect 11518 10911 11574 10920
rect 11028 10906 11034 10908
rect 11090 10906 11114 10908
rect 11170 10906 11194 10908
rect 11250 10906 11274 10908
rect 11330 10906 11336 10908
rect 11090 10854 11092 10906
rect 11272 10854 11274 10906
rect 11028 10852 11034 10854
rect 11090 10852 11114 10854
rect 11170 10852 11194 10854
rect 11250 10852 11274 10854
rect 11330 10852 11336 10854
rect 11028 10843 11336 10852
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10244 8566 10272 10134
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10336 9382 10364 9862
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10368 9276 10676 9285
rect 10368 9274 10374 9276
rect 10430 9274 10454 9276
rect 10510 9274 10534 9276
rect 10590 9274 10614 9276
rect 10670 9274 10676 9276
rect 10430 9222 10432 9274
rect 10612 9222 10614 9274
rect 10368 9220 10374 9222
rect 10430 9220 10454 9222
rect 10510 9220 10534 9222
rect 10590 9220 10614 9222
rect 10670 9220 10676 9222
rect 10368 9211 10676 9220
rect 10704 9042 10732 9318
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10796 8922 10824 9930
rect 11028 9820 11336 9829
rect 11028 9818 11034 9820
rect 11090 9818 11114 9820
rect 11170 9818 11194 9820
rect 11250 9818 11274 9820
rect 11330 9818 11336 9820
rect 11090 9766 11092 9818
rect 11272 9766 11274 9818
rect 11028 9764 11034 9766
rect 11090 9764 11114 9766
rect 11170 9764 11194 9766
rect 11250 9764 11274 9766
rect 11330 9764 11336 9766
rect 11028 9755 11336 9764
rect 11532 9625 11560 9998
rect 11624 9926 11652 11698
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11518 9616 11574 9625
rect 11518 9551 11574 9560
rect 10704 8906 10824 8922
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10692 8900 10824 8906
rect 10744 8894 10824 8900
rect 10692 8842 10744 8848
rect 10612 8634 10640 8842
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10704 8498 10732 8842
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10796 8498 10824 8774
rect 10888 8634 10916 8774
rect 11028 8732 11336 8741
rect 11028 8730 11034 8732
rect 11090 8730 11114 8732
rect 11170 8730 11194 8732
rect 11250 8730 11274 8732
rect 11330 8730 11336 8732
rect 11090 8678 11092 8730
rect 11272 8678 11274 8730
rect 11028 8676 11034 8678
rect 11090 8676 11114 8678
rect 11170 8676 11194 8678
rect 11250 8676 11274 8678
rect 11330 8676 11336 8678
rect 11028 8667 11336 8676
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10368 8188 10676 8197
rect 10368 8186 10374 8188
rect 10430 8186 10454 8188
rect 10510 8186 10534 8188
rect 10590 8186 10614 8188
rect 10670 8186 10676 8188
rect 10430 8134 10432 8186
rect 10612 8134 10614 8186
rect 10368 8132 10374 8134
rect 10430 8132 10454 8134
rect 10510 8132 10534 8134
rect 10590 8132 10614 8134
rect 10670 8132 10676 8134
rect 10368 8123 10676 8132
rect 10368 7100 10676 7109
rect 10368 7098 10374 7100
rect 10430 7098 10454 7100
rect 10510 7098 10534 7100
rect 10590 7098 10614 7100
rect 10670 7098 10676 7100
rect 10430 7046 10432 7098
rect 10612 7046 10614 7098
rect 10368 7044 10374 7046
rect 10430 7044 10454 7046
rect 10510 7044 10534 7046
rect 10590 7044 10614 7046
rect 10670 7044 10676 7046
rect 10368 7035 10676 7044
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10414 6896 10470 6905
rect 10244 5846 10272 6870
rect 10414 6831 10470 6840
rect 10428 6798 10456 6831
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 6118 10364 6666
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6254 10456 6598
rect 10520 6322 10548 6938
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10600 6316 10652 6322
rect 10704 6304 10732 8434
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6361 10824 6666
rect 10888 6662 10916 8230
rect 11028 7644 11336 7653
rect 11028 7642 11034 7644
rect 11090 7642 11114 7644
rect 11170 7642 11194 7644
rect 11250 7642 11274 7644
rect 11330 7642 11336 7644
rect 11090 7590 11092 7642
rect 11272 7590 11274 7642
rect 11028 7588 11034 7590
rect 11090 7588 11114 7590
rect 11170 7588 11194 7590
rect 11250 7588 11274 7590
rect 11330 7588 11336 7590
rect 11028 7579 11336 7588
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 6798 11008 7414
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11256 6905 11284 7346
rect 11440 7002 11468 8502
rect 11518 8256 11574 8265
rect 11518 8191 11574 8200
rect 11532 7886 11560 8191
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11242 6896 11298 6905
rect 11242 6831 11298 6840
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 11426 6624 11482 6633
rect 11028 6556 11336 6565
rect 11426 6559 11482 6568
rect 11028 6554 11034 6556
rect 11090 6554 11114 6556
rect 11170 6554 11194 6556
rect 11250 6554 11274 6556
rect 11330 6554 11336 6556
rect 11090 6502 11092 6554
rect 11272 6502 11274 6554
rect 11028 6500 11034 6502
rect 11090 6500 11114 6502
rect 11170 6500 11194 6502
rect 11250 6500 11274 6502
rect 11330 6500 11336 6502
rect 11028 6491 11336 6500
rect 11152 6384 11204 6390
rect 10600 6258 10652 6264
rect 10684 6276 10732 6304
rect 10782 6352 10838 6361
rect 11152 6326 11204 6332
rect 10782 6287 10838 6296
rect 10876 6316 10928 6322
rect 10416 6248 10468 6254
rect 10612 6225 10640 6258
rect 10416 6190 10468 6196
rect 10598 6216 10654 6225
rect 10598 6151 10654 6160
rect 10684 6168 10712 6276
rect 10876 6258 10928 6264
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10782 6216 10838 6225
rect 10684 6140 10732 6168
rect 10782 6151 10838 6160
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10368 6012 10676 6021
rect 10368 6010 10374 6012
rect 10430 6010 10454 6012
rect 10510 6010 10534 6012
rect 10590 6010 10614 6012
rect 10670 6010 10676 6012
rect 10430 5958 10432 6010
rect 10612 5958 10614 6010
rect 10368 5956 10374 5958
rect 10430 5956 10454 5958
rect 10510 5956 10534 5958
rect 10590 5956 10614 5958
rect 10670 5956 10676 5958
rect 10368 5947 10676 5956
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10506 5808 10562 5817
rect 10506 5743 10562 5752
rect 10230 5672 10286 5681
rect 10140 5636 10192 5642
rect 10230 5607 10286 5616
rect 10140 5578 10192 5584
rect 10244 5370 10272 5607
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10520 5234 10548 5743
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10060 4826 10088 5170
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10244 4758 10272 5170
rect 10612 5012 10640 5850
rect 10704 5710 10732 6140
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10796 5574 10824 6151
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10612 4984 10732 5012
rect 10368 4924 10676 4933
rect 10368 4922 10374 4924
rect 10430 4922 10454 4924
rect 10510 4922 10534 4924
rect 10590 4922 10614 4924
rect 10670 4922 10676 4924
rect 10430 4870 10432 4922
rect 10612 4870 10614 4922
rect 10368 4868 10374 4870
rect 10430 4868 10454 4870
rect 10510 4868 10534 4870
rect 10590 4868 10614 4870
rect 10670 4868 10676 4870
rect 10368 4859 10676 4868
rect 10704 4758 10732 4984
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10704 4570 10732 4694
rect 10796 4622 10824 5510
rect 10520 4554 10732 4570
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10508 4548 10732 4554
rect 10560 4542 10732 4548
rect 10508 4490 10560 4496
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10060 3194 10088 4014
rect 10152 3534 10180 4422
rect 10336 4078 10364 4490
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3738 10272 3878
rect 10368 3836 10676 3845
rect 10368 3834 10374 3836
rect 10430 3834 10454 3836
rect 10510 3834 10534 3836
rect 10590 3834 10614 3836
rect 10670 3834 10676 3836
rect 10430 3782 10432 3834
rect 10612 3782 10614 3834
rect 10368 3780 10374 3782
rect 10430 3780 10454 3782
rect 10510 3780 10534 3782
rect 10590 3780 10614 3782
rect 10670 3780 10676 3782
rect 10368 3771 10676 3780
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10704 3602 10732 4422
rect 10796 4214 10824 4558
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10428 3126 10456 3334
rect 10888 3194 10916 6258
rect 11072 6118 11100 6258
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11164 5914 11192 6326
rect 11440 6304 11468 6559
rect 11348 6276 11468 6304
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11348 5710 11376 6276
rect 11532 6236 11560 6734
rect 11440 6208 11560 6236
rect 11336 5704 11388 5710
rect 11334 5672 11336 5681
rect 11388 5672 11390 5681
rect 11334 5607 11390 5616
rect 11028 5468 11336 5477
rect 11028 5466 11034 5468
rect 11090 5466 11114 5468
rect 11170 5466 11194 5468
rect 11250 5466 11274 5468
rect 11330 5466 11336 5468
rect 11090 5414 11092 5466
rect 11272 5414 11274 5466
rect 11028 5412 11034 5414
rect 11090 5412 11114 5414
rect 11170 5412 11194 5414
rect 11250 5412 11274 5414
rect 11330 5412 11336 5414
rect 11028 5403 11336 5412
rect 11440 5386 11468 6208
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11532 5545 11560 5646
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11518 5536 11574 5545
rect 11518 5471 11574 5480
rect 11440 5358 11560 5386
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10980 4706 11008 4966
rect 10980 4678 11100 4706
rect 11072 4622 11100 4678
rect 11256 4622 11284 4966
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11028 4380 11336 4389
rect 11028 4378 11034 4380
rect 11090 4378 11114 4380
rect 11170 4378 11194 4380
rect 11250 4378 11274 4380
rect 11330 4378 11336 4380
rect 11090 4326 11092 4378
rect 11272 4326 11274 4378
rect 11028 4324 11034 4326
rect 11090 4324 11114 4326
rect 11170 4324 11194 4326
rect 11250 4324 11274 4326
rect 11330 4324 11336 4326
rect 11028 4315 11336 4324
rect 11440 4185 11468 5170
rect 11426 4176 11482 4185
rect 11426 4111 11482 4120
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11028 3292 11336 3301
rect 11028 3290 11034 3292
rect 11090 3290 11114 3292
rect 11170 3290 11194 3292
rect 11250 3290 11274 3292
rect 11330 3290 11336 3292
rect 11090 3238 11092 3290
rect 11272 3238 11274 3290
rect 11028 3236 11034 3238
rect 11090 3236 11114 3238
rect 11170 3236 11194 3238
rect 11250 3236 11274 3238
rect 11330 3236 11336 3238
rect 11028 3227 11336 3236
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 10368 2748 10676 2757
rect 10368 2746 10374 2748
rect 10430 2746 10454 2748
rect 10510 2746 10534 2748
rect 10590 2746 10614 2748
rect 10670 2746 10676 2748
rect 10430 2694 10432 2746
rect 10612 2694 10614 2746
rect 10368 2692 10374 2694
rect 10430 2692 10454 2694
rect 10510 2692 10534 2694
rect 10590 2692 10614 2694
rect 10670 2692 10676 2694
rect 10368 2683 10676 2692
rect 10796 2650 10824 2994
rect 11348 2825 11376 2994
rect 11334 2816 11390 2825
rect 11334 2751 11390 2760
rect 11440 2650 11468 3946
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11532 2582 11560 5358
rect 11624 3194 11652 5578
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3804 1550 3924 1578
rect 3896 800 3924 1550
rect 5184 800 5212 2382
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 5646 2204 5954 2213
rect 5646 2202 5652 2204
rect 5708 2202 5732 2204
rect 5788 2202 5812 2204
rect 5868 2202 5892 2204
rect 5948 2202 5954 2204
rect 5708 2150 5710 2202
rect 5890 2150 5892 2202
rect 5646 2148 5652 2150
rect 5708 2148 5732 2150
rect 5788 2148 5812 2150
rect 5868 2148 5892 2150
rect 5948 2148 5954 2150
rect 5646 2139 5954 2148
rect 6472 800 6500 2314
rect 7760 800 7788 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 8337 2204 8645 2213
rect 8337 2202 8343 2204
rect 8399 2202 8423 2204
rect 8479 2202 8503 2204
rect 8559 2202 8583 2204
rect 8639 2202 8645 2204
rect 8399 2150 8401 2202
rect 8581 2150 8583 2202
rect 8337 2148 8343 2150
rect 8399 2148 8423 2150
rect 8479 2148 8503 2150
rect 8559 2148 8583 2150
rect 8639 2148 8645 2150
rect 8337 2139 8645 2148
rect 9048 800 9076 2246
rect 10428 1306 10456 2382
rect 11028 2204 11336 2213
rect 11028 2202 11034 2204
rect 11090 2202 11114 2204
rect 11170 2202 11194 2204
rect 11250 2202 11274 2204
rect 11330 2202 11336 2204
rect 11090 2150 11092 2202
rect 11272 2150 11274 2202
rect 11028 2148 11034 2150
rect 11090 2148 11114 2150
rect 11170 2148 11194 2150
rect 11250 2148 11274 2150
rect 11330 2148 11336 2150
rect 11028 2139 11336 2148
rect 11440 1465 11468 2450
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11426 1456 11482 1465
rect 11426 1391 11482 1400
rect 10336 1278 10456 1306
rect 10336 800 10364 1278
rect 11624 800 11652 2382
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12912 800 12940 2314
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
<< via2 >>
rect 1030 12280 1086 12336
rect 1490 13640 1546 13696
rect 2301 12538 2357 12540
rect 2381 12538 2437 12540
rect 2461 12538 2517 12540
rect 2541 12538 2597 12540
rect 2301 12486 2347 12538
rect 2347 12486 2357 12538
rect 2381 12486 2411 12538
rect 2411 12486 2423 12538
rect 2423 12486 2437 12538
rect 2461 12486 2475 12538
rect 2475 12486 2487 12538
rect 2487 12486 2517 12538
rect 2541 12486 2551 12538
rect 2551 12486 2597 12538
rect 2301 12484 2357 12486
rect 2381 12484 2437 12486
rect 2461 12484 2517 12486
rect 2541 12484 2597 12486
rect 4992 12538 5048 12540
rect 5072 12538 5128 12540
rect 5152 12538 5208 12540
rect 5232 12538 5288 12540
rect 4992 12486 5038 12538
rect 5038 12486 5048 12538
rect 5072 12486 5102 12538
rect 5102 12486 5114 12538
rect 5114 12486 5128 12538
rect 5152 12486 5166 12538
rect 5166 12486 5178 12538
rect 5178 12486 5208 12538
rect 5232 12486 5242 12538
rect 5242 12486 5288 12538
rect 4992 12484 5048 12486
rect 5072 12484 5128 12486
rect 5152 12484 5208 12486
rect 5232 12484 5288 12486
rect 938 10920 994 10976
rect 1398 9560 1454 9616
rect 1858 11636 1860 11656
rect 1860 11636 1912 11656
rect 1912 11636 1914 11656
rect 1858 11600 1914 11636
rect 2301 11450 2357 11452
rect 2381 11450 2437 11452
rect 2461 11450 2517 11452
rect 2541 11450 2597 11452
rect 2301 11398 2347 11450
rect 2347 11398 2357 11450
rect 2381 11398 2411 11450
rect 2411 11398 2423 11450
rect 2423 11398 2437 11450
rect 2461 11398 2475 11450
rect 2475 11398 2487 11450
rect 2487 11398 2517 11450
rect 2541 11398 2551 11450
rect 2551 11398 2597 11450
rect 2301 11396 2357 11398
rect 2381 11396 2437 11398
rect 2461 11396 2517 11398
rect 2541 11396 2597 11398
rect 2961 11994 3017 11996
rect 3041 11994 3097 11996
rect 3121 11994 3177 11996
rect 3201 11994 3257 11996
rect 2961 11942 3007 11994
rect 3007 11942 3017 11994
rect 3041 11942 3071 11994
rect 3071 11942 3083 11994
rect 3083 11942 3097 11994
rect 3121 11942 3135 11994
rect 3135 11942 3147 11994
rect 3147 11942 3177 11994
rect 3201 11942 3211 11994
rect 3211 11942 3257 11994
rect 2961 11940 3017 11942
rect 3041 11940 3097 11942
rect 3121 11940 3177 11942
rect 3201 11940 3257 11942
rect 2961 10906 3017 10908
rect 3041 10906 3097 10908
rect 3121 10906 3177 10908
rect 3201 10906 3257 10908
rect 2961 10854 3007 10906
rect 3007 10854 3017 10906
rect 3041 10854 3071 10906
rect 3071 10854 3083 10906
rect 3083 10854 3097 10906
rect 3121 10854 3135 10906
rect 3135 10854 3147 10906
rect 3147 10854 3177 10906
rect 3201 10854 3211 10906
rect 3211 10854 3257 10906
rect 2961 10852 3017 10854
rect 3041 10852 3097 10854
rect 3121 10852 3177 10854
rect 3201 10852 3257 10854
rect 2301 10362 2357 10364
rect 2381 10362 2437 10364
rect 2461 10362 2517 10364
rect 2541 10362 2597 10364
rect 2301 10310 2347 10362
rect 2347 10310 2357 10362
rect 2381 10310 2411 10362
rect 2411 10310 2423 10362
rect 2423 10310 2437 10362
rect 2461 10310 2475 10362
rect 2475 10310 2487 10362
rect 2487 10310 2517 10362
rect 2541 10310 2551 10362
rect 2551 10310 2597 10362
rect 2301 10308 2357 10310
rect 2381 10308 2437 10310
rect 2461 10308 2517 10310
rect 2541 10308 2597 10310
rect 1398 8200 1454 8256
rect 1398 6840 1454 6896
rect 938 5480 994 5536
rect 1306 4120 1362 4176
rect 938 2760 994 2816
rect 2961 9818 3017 9820
rect 3041 9818 3097 9820
rect 3121 9818 3177 9820
rect 3201 9818 3257 9820
rect 2961 9766 3007 9818
rect 3007 9766 3017 9818
rect 3041 9766 3071 9818
rect 3071 9766 3083 9818
rect 3083 9766 3097 9818
rect 3121 9766 3135 9818
rect 3135 9766 3147 9818
rect 3147 9766 3177 9818
rect 3201 9766 3211 9818
rect 3211 9766 3257 9818
rect 2961 9764 3017 9766
rect 3041 9764 3097 9766
rect 3121 9764 3177 9766
rect 3201 9764 3257 9766
rect 2301 9274 2357 9276
rect 2381 9274 2437 9276
rect 2461 9274 2517 9276
rect 2541 9274 2597 9276
rect 2301 9222 2347 9274
rect 2347 9222 2357 9274
rect 2381 9222 2411 9274
rect 2411 9222 2423 9274
rect 2423 9222 2437 9274
rect 2461 9222 2475 9274
rect 2475 9222 2487 9274
rect 2487 9222 2517 9274
rect 2541 9222 2551 9274
rect 2551 9222 2597 9274
rect 2301 9220 2357 9222
rect 2381 9220 2437 9222
rect 2461 9220 2517 9222
rect 2541 9220 2597 9222
rect 1674 5208 1730 5264
rect 1582 4004 1638 4040
rect 1582 3984 1584 4004
rect 1584 3984 1636 4004
rect 1636 3984 1638 4004
rect 2301 8186 2357 8188
rect 2381 8186 2437 8188
rect 2461 8186 2517 8188
rect 2541 8186 2597 8188
rect 2301 8134 2347 8186
rect 2347 8134 2357 8186
rect 2381 8134 2411 8186
rect 2411 8134 2423 8186
rect 2423 8134 2437 8186
rect 2461 8134 2475 8186
rect 2475 8134 2487 8186
rect 2487 8134 2517 8186
rect 2541 8134 2551 8186
rect 2551 8134 2597 8186
rect 2301 8132 2357 8134
rect 2381 8132 2437 8134
rect 2461 8132 2517 8134
rect 2541 8132 2597 8134
rect 2961 8730 3017 8732
rect 3041 8730 3097 8732
rect 3121 8730 3177 8732
rect 3201 8730 3257 8732
rect 2961 8678 3007 8730
rect 3007 8678 3017 8730
rect 3041 8678 3071 8730
rect 3071 8678 3083 8730
rect 3083 8678 3097 8730
rect 3121 8678 3135 8730
rect 3135 8678 3147 8730
rect 3147 8678 3177 8730
rect 3201 8678 3211 8730
rect 3211 8678 3257 8730
rect 2961 8676 3017 8678
rect 3041 8676 3097 8678
rect 3121 8676 3177 8678
rect 3201 8676 3257 8678
rect 3238 7964 3240 7984
rect 3240 7964 3292 7984
rect 3292 7964 3294 7984
rect 3238 7928 3294 7964
rect 2961 7642 3017 7644
rect 3041 7642 3097 7644
rect 3121 7642 3177 7644
rect 3201 7642 3257 7644
rect 2961 7590 3007 7642
rect 3007 7590 3017 7642
rect 3041 7590 3071 7642
rect 3071 7590 3083 7642
rect 3083 7590 3097 7642
rect 3121 7590 3135 7642
rect 3135 7590 3147 7642
rect 3147 7590 3177 7642
rect 3201 7590 3211 7642
rect 3211 7590 3257 7642
rect 2961 7588 3017 7590
rect 3041 7588 3097 7590
rect 3121 7588 3177 7590
rect 3201 7588 3257 7590
rect 3514 7792 3570 7848
rect 2301 7098 2357 7100
rect 2381 7098 2437 7100
rect 2461 7098 2517 7100
rect 2541 7098 2597 7100
rect 2301 7046 2347 7098
rect 2347 7046 2357 7098
rect 2381 7046 2411 7098
rect 2411 7046 2423 7098
rect 2423 7046 2437 7098
rect 2461 7046 2475 7098
rect 2475 7046 2487 7098
rect 2487 7046 2517 7098
rect 2541 7046 2551 7098
rect 2551 7046 2597 7098
rect 2301 7044 2357 7046
rect 2381 7044 2437 7046
rect 2461 7044 2517 7046
rect 2541 7044 2597 7046
rect 2301 6010 2357 6012
rect 2381 6010 2437 6012
rect 2461 6010 2517 6012
rect 2541 6010 2597 6012
rect 2301 5958 2347 6010
rect 2347 5958 2357 6010
rect 2381 5958 2411 6010
rect 2411 5958 2423 6010
rect 2423 5958 2437 6010
rect 2461 5958 2475 6010
rect 2475 5958 2487 6010
rect 2487 5958 2517 6010
rect 2541 5958 2551 6010
rect 2551 5958 2597 6010
rect 2301 5956 2357 5958
rect 2381 5956 2437 5958
rect 2461 5956 2517 5958
rect 2541 5956 2597 5958
rect 2301 4922 2357 4924
rect 2381 4922 2437 4924
rect 2461 4922 2517 4924
rect 2541 4922 2597 4924
rect 2301 4870 2347 4922
rect 2347 4870 2357 4922
rect 2381 4870 2411 4922
rect 2411 4870 2423 4922
rect 2423 4870 2437 4922
rect 2461 4870 2475 4922
rect 2475 4870 2487 4922
rect 2487 4870 2517 4922
rect 2541 4870 2551 4922
rect 2551 4870 2597 4922
rect 2301 4868 2357 4870
rect 2381 4868 2437 4870
rect 2461 4868 2517 4870
rect 2541 4868 2597 4870
rect 2301 3834 2357 3836
rect 2381 3834 2437 3836
rect 2461 3834 2517 3836
rect 2541 3834 2597 3836
rect 2301 3782 2347 3834
rect 2347 3782 2357 3834
rect 2381 3782 2411 3834
rect 2411 3782 2423 3834
rect 2423 3782 2437 3834
rect 2461 3782 2475 3834
rect 2475 3782 2487 3834
rect 2487 3782 2517 3834
rect 2541 3782 2551 3834
rect 2551 3782 2597 3834
rect 2301 3780 2357 3782
rect 2381 3780 2437 3782
rect 2461 3780 2517 3782
rect 2541 3780 2597 3782
rect 2594 3032 2650 3088
rect 2318 2916 2374 2952
rect 2318 2896 2320 2916
rect 2320 2896 2372 2916
rect 2372 2896 2374 2916
rect 2301 2746 2357 2748
rect 2381 2746 2437 2748
rect 2461 2746 2517 2748
rect 2541 2746 2597 2748
rect 2301 2694 2347 2746
rect 2347 2694 2357 2746
rect 2381 2694 2411 2746
rect 2411 2694 2423 2746
rect 2423 2694 2437 2746
rect 2461 2694 2475 2746
rect 2475 2694 2487 2746
rect 2487 2694 2517 2746
rect 2541 2694 2551 2746
rect 2551 2694 2597 2746
rect 2301 2692 2357 2694
rect 2381 2692 2437 2694
rect 2461 2692 2517 2694
rect 2541 2692 2597 2694
rect 2961 6554 3017 6556
rect 3041 6554 3097 6556
rect 3121 6554 3177 6556
rect 3201 6554 3257 6556
rect 2961 6502 3007 6554
rect 3007 6502 3017 6554
rect 3041 6502 3071 6554
rect 3071 6502 3083 6554
rect 3083 6502 3097 6554
rect 3121 6502 3135 6554
rect 3135 6502 3147 6554
rect 3147 6502 3177 6554
rect 3201 6502 3211 6554
rect 3211 6502 3257 6554
rect 2961 6500 3017 6502
rect 3041 6500 3097 6502
rect 3121 6500 3177 6502
rect 3201 6500 3257 6502
rect 4250 11076 4306 11112
rect 4250 11056 4252 11076
rect 4252 11056 4304 11076
rect 4304 11056 4306 11076
rect 3606 6160 3662 6216
rect 2961 5466 3017 5468
rect 3041 5466 3097 5468
rect 3121 5466 3177 5468
rect 3201 5466 3257 5468
rect 2961 5414 3007 5466
rect 3007 5414 3017 5466
rect 3041 5414 3071 5466
rect 3071 5414 3083 5466
rect 3083 5414 3097 5466
rect 3121 5414 3135 5466
rect 3135 5414 3147 5466
rect 3147 5414 3177 5466
rect 3201 5414 3211 5466
rect 3211 5414 3257 5466
rect 2961 5412 3017 5414
rect 3041 5412 3097 5414
rect 3121 5412 3177 5414
rect 3201 5412 3257 5414
rect 3330 4528 3386 4584
rect 2961 4378 3017 4380
rect 3041 4378 3097 4380
rect 3121 4378 3177 4380
rect 3201 4378 3257 4380
rect 2961 4326 3007 4378
rect 3007 4326 3017 4378
rect 3041 4326 3071 4378
rect 3071 4326 3083 4378
rect 3083 4326 3097 4378
rect 3121 4326 3135 4378
rect 3135 4326 3147 4378
rect 3147 4326 3177 4378
rect 3201 4326 3211 4378
rect 3211 4326 3257 4378
rect 2961 4324 3017 4326
rect 3041 4324 3097 4326
rect 3121 4324 3177 4326
rect 3201 4324 3257 4326
rect 2961 3290 3017 3292
rect 3041 3290 3097 3292
rect 3121 3290 3177 3292
rect 3201 3290 3257 3292
rect 2961 3238 3007 3290
rect 3007 3238 3017 3290
rect 3041 3238 3071 3290
rect 3071 3238 3083 3290
rect 3083 3238 3097 3290
rect 3121 3238 3135 3290
rect 3135 3238 3147 3290
rect 3147 3238 3177 3290
rect 3201 3238 3211 3290
rect 3211 3238 3257 3290
rect 2961 3236 3017 3238
rect 3041 3236 3097 3238
rect 3121 3236 3177 3238
rect 3201 3236 3257 3238
rect 4618 7928 4674 7984
rect 4992 11450 5048 11452
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 4992 11398 5038 11450
rect 5038 11398 5048 11450
rect 5072 11398 5102 11450
rect 5102 11398 5114 11450
rect 5114 11398 5128 11450
rect 5152 11398 5166 11450
rect 5166 11398 5178 11450
rect 5178 11398 5208 11450
rect 5232 11398 5242 11450
rect 5242 11398 5288 11450
rect 4992 11396 5048 11398
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 4992 10362 5048 10364
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 4992 10310 5038 10362
rect 5038 10310 5048 10362
rect 5072 10310 5102 10362
rect 5102 10310 5114 10362
rect 5114 10310 5128 10362
rect 5152 10310 5166 10362
rect 5166 10310 5178 10362
rect 5178 10310 5208 10362
rect 5232 10310 5242 10362
rect 5242 10310 5288 10362
rect 4992 10308 5048 10310
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 4992 9274 5048 9276
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 4992 9222 5038 9274
rect 5038 9222 5048 9274
rect 5072 9222 5102 9274
rect 5102 9222 5114 9274
rect 5114 9222 5128 9274
rect 5152 9222 5166 9274
rect 5166 9222 5178 9274
rect 5178 9222 5208 9274
rect 5232 9222 5242 9274
rect 5242 9222 5288 9274
rect 4992 9220 5048 9222
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 7683 12538 7739 12540
rect 7763 12538 7819 12540
rect 7843 12538 7899 12540
rect 7923 12538 7979 12540
rect 7683 12486 7729 12538
rect 7729 12486 7739 12538
rect 7763 12486 7793 12538
rect 7793 12486 7805 12538
rect 7805 12486 7819 12538
rect 7843 12486 7857 12538
rect 7857 12486 7869 12538
rect 7869 12486 7899 12538
rect 7923 12486 7933 12538
rect 7933 12486 7979 12538
rect 7683 12484 7739 12486
rect 7763 12484 7819 12486
rect 7843 12484 7899 12486
rect 7923 12484 7979 12486
rect 5652 11994 5708 11996
rect 5732 11994 5788 11996
rect 5812 11994 5868 11996
rect 5892 11994 5948 11996
rect 5652 11942 5698 11994
rect 5698 11942 5708 11994
rect 5732 11942 5762 11994
rect 5762 11942 5774 11994
rect 5774 11942 5788 11994
rect 5812 11942 5826 11994
rect 5826 11942 5838 11994
rect 5838 11942 5868 11994
rect 5892 11942 5902 11994
rect 5902 11942 5948 11994
rect 5652 11940 5708 11942
rect 5732 11940 5788 11942
rect 5812 11940 5868 11942
rect 5892 11940 5948 11942
rect 5652 10906 5708 10908
rect 5732 10906 5788 10908
rect 5812 10906 5868 10908
rect 5892 10906 5948 10908
rect 5652 10854 5698 10906
rect 5698 10854 5708 10906
rect 5732 10854 5762 10906
rect 5762 10854 5774 10906
rect 5774 10854 5788 10906
rect 5812 10854 5826 10906
rect 5826 10854 5838 10906
rect 5838 10854 5868 10906
rect 5892 10854 5902 10906
rect 5902 10854 5948 10906
rect 5652 10852 5708 10854
rect 5732 10852 5788 10854
rect 5812 10852 5868 10854
rect 5892 10852 5948 10854
rect 5652 9818 5708 9820
rect 5732 9818 5788 9820
rect 5812 9818 5868 9820
rect 5892 9818 5948 9820
rect 5652 9766 5698 9818
rect 5698 9766 5708 9818
rect 5732 9766 5762 9818
rect 5762 9766 5774 9818
rect 5774 9766 5788 9818
rect 5812 9766 5826 9818
rect 5826 9766 5838 9818
rect 5838 9766 5868 9818
rect 5892 9766 5902 9818
rect 5902 9766 5948 9818
rect 5652 9764 5708 9766
rect 5732 9764 5788 9766
rect 5812 9764 5868 9766
rect 5892 9764 5948 9766
rect 5170 8336 5226 8392
rect 4992 8186 5048 8188
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 4992 8134 5038 8186
rect 5038 8134 5048 8186
rect 5072 8134 5102 8186
rect 5102 8134 5114 8186
rect 5114 8134 5128 8186
rect 5152 8134 5166 8186
rect 5166 8134 5178 8186
rect 5178 8134 5208 8186
rect 5232 8134 5242 8186
rect 5242 8134 5288 8186
rect 4992 8132 5048 8134
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 4250 3476 4252 3496
rect 4252 3476 4304 3496
rect 4304 3476 4306 3496
rect 4250 3440 4306 3476
rect 2961 2202 3017 2204
rect 3041 2202 3097 2204
rect 3121 2202 3177 2204
rect 3201 2202 3257 2204
rect 2961 2150 3007 2202
rect 3007 2150 3017 2202
rect 3041 2150 3071 2202
rect 3071 2150 3083 2202
rect 3083 2150 3097 2202
rect 3121 2150 3135 2202
rect 3135 2150 3147 2202
rect 3147 2150 3177 2202
rect 3201 2150 3211 2202
rect 3211 2150 3257 2202
rect 2961 2148 3017 2150
rect 3041 2148 3097 2150
rect 3121 2148 3177 2150
rect 3201 2148 3257 2150
rect 1398 1400 1454 1456
rect 4992 7098 5048 7100
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 4992 7046 5038 7098
rect 5038 7046 5048 7098
rect 5072 7046 5102 7098
rect 5102 7046 5114 7098
rect 5114 7046 5128 7098
rect 5152 7046 5166 7098
rect 5166 7046 5178 7098
rect 5178 7046 5208 7098
rect 5232 7046 5242 7098
rect 5242 7046 5288 7098
rect 4992 7044 5048 7046
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 6458 11600 6514 11656
rect 6366 8880 6422 8936
rect 5652 8730 5708 8732
rect 5732 8730 5788 8732
rect 5812 8730 5868 8732
rect 5892 8730 5948 8732
rect 5652 8678 5698 8730
rect 5698 8678 5708 8730
rect 5732 8678 5762 8730
rect 5762 8678 5774 8730
rect 5774 8678 5788 8730
rect 5812 8678 5826 8730
rect 5826 8678 5838 8730
rect 5838 8678 5868 8730
rect 5892 8678 5902 8730
rect 5902 8678 5948 8730
rect 5652 8676 5708 8678
rect 5732 8676 5788 8678
rect 5812 8676 5868 8678
rect 5892 8676 5948 8678
rect 5652 7642 5708 7644
rect 5732 7642 5788 7644
rect 5812 7642 5868 7644
rect 5892 7642 5948 7644
rect 5652 7590 5698 7642
rect 5698 7590 5708 7642
rect 5732 7590 5762 7642
rect 5762 7590 5774 7642
rect 5774 7590 5788 7642
rect 5812 7590 5826 7642
rect 5826 7590 5838 7642
rect 5838 7590 5868 7642
rect 5892 7590 5902 7642
rect 5902 7590 5948 7642
rect 5652 7588 5708 7590
rect 5732 7588 5788 7590
rect 5812 7588 5868 7590
rect 5892 7588 5948 7590
rect 4992 6010 5048 6012
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 4992 5958 5038 6010
rect 5038 5958 5048 6010
rect 5072 5958 5102 6010
rect 5102 5958 5114 6010
rect 5114 5958 5128 6010
rect 5152 5958 5166 6010
rect 5166 5958 5178 6010
rect 5178 5958 5208 6010
rect 5232 5958 5242 6010
rect 5242 5958 5288 6010
rect 4992 5956 5048 5958
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 5652 6554 5708 6556
rect 5732 6554 5788 6556
rect 5812 6554 5868 6556
rect 5892 6554 5948 6556
rect 5652 6502 5698 6554
rect 5698 6502 5708 6554
rect 5732 6502 5762 6554
rect 5762 6502 5774 6554
rect 5774 6502 5788 6554
rect 5812 6502 5826 6554
rect 5826 6502 5838 6554
rect 5838 6502 5868 6554
rect 5892 6502 5902 6554
rect 5902 6502 5948 6554
rect 5652 6500 5708 6502
rect 5732 6500 5788 6502
rect 5812 6500 5868 6502
rect 5892 6500 5948 6502
rect 5630 6024 5686 6080
rect 5446 5244 5448 5264
rect 5448 5244 5500 5264
rect 5500 5244 5502 5264
rect 5446 5208 5502 5244
rect 5652 5466 5708 5468
rect 5732 5466 5788 5468
rect 5812 5466 5868 5468
rect 5892 5466 5948 5468
rect 5652 5414 5698 5466
rect 5698 5414 5708 5466
rect 5732 5414 5762 5466
rect 5762 5414 5774 5466
rect 5774 5414 5788 5466
rect 5812 5414 5826 5466
rect 5826 5414 5838 5466
rect 5838 5414 5868 5466
rect 5892 5414 5902 5466
rect 5902 5414 5948 5466
rect 5652 5412 5708 5414
rect 5732 5412 5788 5414
rect 5812 5412 5868 5414
rect 5892 5412 5948 5414
rect 4992 4922 5048 4924
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 4992 4870 5038 4922
rect 5038 4870 5048 4922
rect 5072 4870 5102 4922
rect 5102 4870 5114 4922
rect 5114 4870 5128 4922
rect 5152 4870 5166 4922
rect 5166 4870 5178 4922
rect 5178 4870 5208 4922
rect 5232 4870 5242 4922
rect 5242 4870 5288 4922
rect 4992 4868 5048 4870
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 4992 3834 5048 3836
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 4992 3782 5038 3834
rect 5038 3782 5048 3834
rect 5072 3782 5102 3834
rect 5102 3782 5114 3834
rect 5114 3782 5128 3834
rect 5152 3782 5166 3834
rect 5166 3782 5178 3834
rect 5178 3782 5208 3834
rect 5232 3782 5242 3834
rect 5242 3782 5288 3834
rect 4992 3780 5048 3782
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5814 4664 5870 4720
rect 5652 4378 5708 4380
rect 5732 4378 5788 4380
rect 5812 4378 5868 4380
rect 5892 4378 5948 4380
rect 5652 4326 5698 4378
rect 5698 4326 5708 4378
rect 5732 4326 5762 4378
rect 5762 4326 5774 4378
rect 5774 4326 5788 4378
rect 5812 4326 5826 4378
rect 5826 4326 5838 4378
rect 5838 4326 5868 4378
rect 5892 4326 5902 4378
rect 5902 4326 5948 4378
rect 5652 4324 5708 4326
rect 5732 4324 5788 4326
rect 5812 4324 5868 4326
rect 5892 4324 5948 4326
rect 5652 3290 5708 3292
rect 5732 3290 5788 3292
rect 5812 3290 5868 3292
rect 5892 3290 5948 3292
rect 5652 3238 5698 3290
rect 5698 3238 5708 3290
rect 5732 3238 5762 3290
rect 5762 3238 5774 3290
rect 5774 3238 5788 3290
rect 5812 3238 5826 3290
rect 5826 3238 5838 3290
rect 5838 3238 5868 3290
rect 5892 3238 5902 3290
rect 5902 3238 5948 3290
rect 5652 3236 5708 3238
rect 5732 3236 5788 3238
rect 5812 3236 5868 3238
rect 5892 3236 5948 3238
rect 6734 8336 6790 8392
rect 11426 13640 11482 13696
rect 8343 11994 8399 11996
rect 8423 11994 8479 11996
rect 8503 11994 8559 11996
rect 8583 11994 8639 11996
rect 8343 11942 8389 11994
rect 8389 11942 8399 11994
rect 8423 11942 8453 11994
rect 8453 11942 8465 11994
rect 8465 11942 8479 11994
rect 8503 11942 8517 11994
rect 8517 11942 8529 11994
rect 8529 11942 8559 11994
rect 8583 11942 8593 11994
rect 8593 11942 8639 11994
rect 8343 11940 8399 11942
rect 8423 11940 8479 11942
rect 8503 11940 8559 11942
rect 8583 11940 8639 11942
rect 6366 5208 6422 5264
rect 6182 4528 6238 4584
rect 6274 3984 6330 4040
rect 6182 3848 6238 3904
rect 5814 3052 5870 3088
rect 5814 3032 5816 3052
rect 5816 3032 5868 3052
rect 5868 3032 5870 3052
rect 4992 2746 5048 2748
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 4992 2694 5038 2746
rect 5038 2694 5048 2746
rect 5072 2694 5102 2746
rect 5102 2694 5114 2746
rect 5114 2694 5128 2746
rect 5152 2694 5166 2746
rect 5166 2694 5178 2746
rect 5178 2694 5208 2746
rect 5232 2694 5242 2746
rect 5242 2694 5288 2746
rect 4992 2692 5048 2694
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 5906 2896 5962 2952
rect 6734 6024 6790 6080
rect 6458 3304 6514 3360
rect 6366 2896 6422 2952
rect 6734 3576 6790 3632
rect 7683 11450 7739 11452
rect 7763 11450 7819 11452
rect 7843 11450 7899 11452
rect 7923 11450 7979 11452
rect 7683 11398 7729 11450
rect 7729 11398 7739 11450
rect 7763 11398 7793 11450
rect 7793 11398 7805 11450
rect 7805 11398 7819 11450
rect 7843 11398 7857 11450
rect 7857 11398 7869 11450
rect 7869 11398 7899 11450
rect 7923 11398 7933 11450
rect 7933 11398 7979 11450
rect 7683 11396 7739 11398
rect 7763 11396 7819 11398
rect 7843 11396 7899 11398
rect 7923 11396 7979 11398
rect 8343 10906 8399 10908
rect 8423 10906 8479 10908
rect 8503 10906 8559 10908
rect 8583 10906 8639 10908
rect 8343 10854 8389 10906
rect 8389 10854 8399 10906
rect 8423 10854 8453 10906
rect 8453 10854 8465 10906
rect 8465 10854 8479 10906
rect 8503 10854 8517 10906
rect 8517 10854 8529 10906
rect 8529 10854 8559 10906
rect 8583 10854 8593 10906
rect 8593 10854 8639 10906
rect 8343 10852 8399 10854
rect 8423 10852 8479 10854
rect 8503 10852 8559 10854
rect 8583 10852 8639 10854
rect 8942 11056 8998 11112
rect 7683 10362 7739 10364
rect 7763 10362 7819 10364
rect 7843 10362 7899 10364
rect 7923 10362 7979 10364
rect 7683 10310 7729 10362
rect 7729 10310 7739 10362
rect 7763 10310 7793 10362
rect 7793 10310 7805 10362
rect 7805 10310 7819 10362
rect 7843 10310 7857 10362
rect 7857 10310 7869 10362
rect 7869 10310 7899 10362
rect 7923 10310 7933 10362
rect 7933 10310 7979 10362
rect 7683 10308 7739 10310
rect 7763 10308 7819 10310
rect 7843 10308 7899 10310
rect 7923 10308 7979 10310
rect 7470 9832 7526 9888
rect 7683 9274 7739 9276
rect 7763 9274 7819 9276
rect 7843 9274 7899 9276
rect 7923 9274 7979 9276
rect 7683 9222 7729 9274
rect 7729 9222 7739 9274
rect 7763 9222 7793 9274
rect 7793 9222 7805 9274
rect 7805 9222 7819 9274
rect 7843 9222 7857 9274
rect 7857 9222 7869 9274
rect 7869 9222 7899 9274
rect 7923 9222 7933 9274
rect 7933 9222 7979 9274
rect 7683 9220 7739 9222
rect 7763 9220 7819 9222
rect 7843 9220 7899 9222
rect 7923 9220 7979 9222
rect 7683 8186 7739 8188
rect 7763 8186 7819 8188
rect 7843 8186 7899 8188
rect 7923 8186 7979 8188
rect 7683 8134 7729 8186
rect 7729 8134 7739 8186
rect 7763 8134 7793 8186
rect 7793 8134 7805 8186
rect 7805 8134 7819 8186
rect 7843 8134 7857 8186
rect 7857 8134 7869 8186
rect 7869 8134 7899 8186
rect 7923 8134 7933 8186
rect 7933 8134 7979 8186
rect 7683 8132 7739 8134
rect 7763 8132 7819 8134
rect 7843 8132 7899 8134
rect 7923 8132 7979 8134
rect 7683 7098 7739 7100
rect 7763 7098 7819 7100
rect 7843 7098 7899 7100
rect 7923 7098 7979 7100
rect 7683 7046 7729 7098
rect 7729 7046 7739 7098
rect 7763 7046 7793 7098
rect 7793 7046 7805 7098
rect 7805 7046 7819 7098
rect 7843 7046 7857 7098
rect 7857 7046 7869 7098
rect 7869 7046 7899 7098
rect 7923 7046 7933 7098
rect 7933 7046 7979 7098
rect 7683 7044 7739 7046
rect 7763 7044 7819 7046
rect 7843 7044 7899 7046
rect 7923 7044 7979 7046
rect 7102 6316 7158 6352
rect 7102 6296 7104 6316
rect 7104 6296 7156 6316
rect 7156 6296 7158 6316
rect 6918 4664 6974 4720
rect 7286 5228 7342 5264
rect 7286 5208 7288 5228
rect 7288 5208 7340 5228
rect 7340 5208 7342 5228
rect 6826 3440 6882 3496
rect 7654 6180 7710 6216
rect 7654 6160 7656 6180
rect 7656 6160 7708 6180
rect 7708 6160 7710 6180
rect 7683 6010 7739 6012
rect 7763 6010 7819 6012
rect 7843 6010 7899 6012
rect 7923 6010 7979 6012
rect 7683 5958 7729 6010
rect 7729 5958 7739 6010
rect 7763 5958 7793 6010
rect 7793 5958 7805 6010
rect 7805 5958 7819 6010
rect 7843 5958 7857 6010
rect 7857 5958 7869 6010
rect 7869 5958 7899 6010
rect 7923 5958 7933 6010
rect 7933 5958 7979 6010
rect 7683 5956 7739 5958
rect 7763 5956 7819 5958
rect 7843 5956 7899 5958
rect 7923 5956 7979 5958
rect 7683 4922 7739 4924
rect 7763 4922 7819 4924
rect 7843 4922 7899 4924
rect 7923 4922 7979 4924
rect 7683 4870 7729 4922
rect 7729 4870 7739 4922
rect 7763 4870 7793 4922
rect 7793 4870 7805 4922
rect 7805 4870 7819 4922
rect 7843 4870 7857 4922
rect 7857 4870 7869 4922
rect 7869 4870 7899 4922
rect 7923 4870 7933 4922
rect 7933 4870 7979 4922
rect 7683 4868 7739 4870
rect 7763 4868 7819 4870
rect 7843 4868 7899 4870
rect 7923 4868 7979 4870
rect 7838 4664 7894 4720
rect 8343 9818 8399 9820
rect 8423 9818 8479 9820
rect 8503 9818 8559 9820
rect 8583 9818 8639 9820
rect 8343 9766 8389 9818
rect 8389 9766 8399 9818
rect 8423 9766 8453 9818
rect 8453 9766 8465 9818
rect 8465 9766 8479 9818
rect 8503 9766 8517 9818
rect 8517 9766 8529 9818
rect 8529 9766 8559 9818
rect 8583 9766 8593 9818
rect 8593 9766 8639 9818
rect 8343 9764 8399 9766
rect 8423 9764 8479 9766
rect 8503 9764 8559 9766
rect 8583 9764 8639 9766
rect 8022 4664 8078 4720
rect 8343 8730 8399 8732
rect 8423 8730 8479 8732
rect 8503 8730 8559 8732
rect 8583 8730 8639 8732
rect 8343 8678 8389 8730
rect 8389 8678 8399 8730
rect 8423 8678 8453 8730
rect 8453 8678 8465 8730
rect 8465 8678 8479 8730
rect 8503 8678 8517 8730
rect 8517 8678 8529 8730
rect 8529 8678 8559 8730
rect 8583 8678 8593 8730
rect 8593 8678 8639 8730
rect 8343 8676 8399 8678
rect 8423 8676 8479 8678
rect 8503 8676 8559 8678
rect 8583 8676 8639 8678
rect 8942 8200 8998 8256
rect 8343 7642 8399 7644
rect 8423 7642 8479 7644
rect 8503 7642 8559 7644
rect 8583 7642 8639 7644
rect 8343 7590 8389 7642
rect 8389 7590 8399 7642
rect 8423 7590 8453 7642
rect 8453 7590 8465 7642
rect 8465 7590 8479 7642
rect 8503 7590 8517 7642
rect 8517 7590 8529 7642
rect 8529 7590 8559 7642
rect 8583 7590 8593 7642
rect 8593 7590 8639 7642
rect 8343 7588 8399 7590
rect 8423 7588 8479 7590
rect 8503 7588 8559 7590
rect 8583 7588 8639 7590
rect 8343 6554 8399 6556
rect 8423 6554 8479 6556
rect 8503 6554 8559 6556
rect 8583 6554 8639 6556
rect 8343 6502 8389 6554
rect 8389 6502 8399 6554
rect 8423 6502 8453 6554
rect 8453 6502 8465 6554
rect 8465 6502 8479 6554
rect 8503 6502 8517 6554
rect 8517 6502 8529 6554
rect 8529 6502 8559 6554
rect 8583 6502 8593 6554
rect 8593 6502 8639 6554
rect 8343 6500 8399 6502
rect 8423 6500 8479 6502
rect 8503 6500 8559 6502
rect 8583 6500 8639 6502
rect 8298 6316 8354 6352
rect 8298 6296 8300 6316
rect 8300 6296 8352 6316
rect 8352 6296 8354 6316
rect 8343 5466 8399 5468
rect 8423 5466 8479 5468
rect 8503 5466 8559 5468
rect 8583 5466 8639 5468
rect 8343 5414 8389 5466
rect 8389 5414 8399 5466
rect 8423 5414 8453 5466
rect 8453 5414 8465 5466
rect 8465 5414 8479 5466
rect 8503 5414 8517 5466
rect 8517 5414 8529 5466
rect 8529 5414 8559 5466
rect 8583 5414 8593 5466
rect 8593 5414 8639 5466
rect 8343 5412 8399 5414
rect 8423 5412 8479 5414
rect 8503 5412 8559 5414
rect 8583 5412 8639 5414
rect 8574 5228 8630 5264
rect 8574 5208 8576 5228
rect 8576 5208 8628 5228
rect 8628 5208 8630 5228
rect 8343 4378 8399 4380
rect 8423 4378 8479 4380
rect 8503 4378 8559 4380
rect 8583 4378 8639 4380
rect 8343 4326 8389 4378
rect 8389 4326 8399 4378
rect 8423 4326 8453 4378
rect 8453 4326 8465 4378
rect 8465 4326 8479 4378
rect 8503 4326 8517 4378
rect 8517 4326 8529 4378
rect 8529 4326 8559 4378
rect 8583 4326 8593 4378
rect 8593 4326 8639 4378
rect 8343 4324 8399 4326
rect 8423 4324 8479 4326
rect 8503 4324 8559 4326
rect 8583 4324 8639 4326
rect 7683 3834 7739 3836
rect 7763 3834 7819 3836
rect 7843 3834 7899 3836
rect 7923 3834 7979 3836
rect 7683 3782 7729 3834
rect 7729 3782 7739 3834
rect 7763 3782 7793 3834
rect 7793 3782 7805 3834
rect 7805 3782 7819 3834
rect 7843 3782 7857 3834
rect 7857 3782 7869 3834
rect 7869 3782 7899 3834
rect 7923 3782 7933 3834
rect 7933 3782 7979 3834
rect 7683 3780 7739 3782
rect 7763 3780 7819 3782
rect 7843 3780 7899 3782
rect 7923 3780 7979 3782
rect 7102 3576 7158 3632
rect 7378 3304 7434 3360
rect 8343 3290 8399 3292
rect 8423 3290 8479 3292
rect 8503 3290 8559 3292
rect 8583 3290 8639 3292
rect 8343 3238 8389 3290
rect 8389 3238 8399 3290
rect 8423 3238 8453 3290
rect 8453 3238 8465 3290
rect 8465 3238 8479 3290
rect 8503 3238 8517 3290
rect 8517 3238 8529 3290
rect 8529 3238 8559 3290
rect 8583 3238 8593 3290
rect 8593 3238 8639 3290
rect 8343 3236 8399 3238
rect 8423 3236 8479 3238
rect 8503 3236 8559 3238
rect 8583 3236 8639 3238
rect 9402 8200 9458 8256
rect 10374 12538 10430 12540
rect 10454 12538 10510 12540
rect 10534 12538 10590 12540
rect 10614 12538 10670 12540
rect 10374 12486 10420 12538
rect 10420 12486 10430 12538
rect 10454 12486 10484 12538
rect 10484 12486 10496 12538
rect 10496 12486 10510 12538
rect 10534 12486 10548 12538
rect 10548 12486 10560 12538
rect 10560 12486 10590 12538
rect 10614 12486 10624 12538
rect 10624 12486 10670 12538
rect 10374 12484 10430 12486
rect 10454 12484 10510 12486
rect 10534 12484 10590 12486
rect 10614 12484 10670 12486
rect 11034 11994 11090 11996
rect 11114 11994 11170 11996
rect 11194 11994 11250 11996
rect 11274 11994 11330 11996
rect 11034 11942 11080 11994
rect 11080 11942 11090 11994
rect 11114 11942 11144 11994
rect 11144 11942 11156 11994
rect 11156 11942 11170 11994
rect 11194 11942 11208 11994
rect 11208 11942 11220 11994
rect 11220 11942 11250 11994
rect 11274 11942 11284 11994
rect 11284 11942 11330 11994
rect 11034 11940 11090 11942
rect 11114 11940 11170 11942
rect 11194 11940 11250 11942
rect 11274 11940 11330 11942
rect 11518 12280 11574 12336
rect 10374 11450 10430 11452
rect 10454 11450 10510 11452
rect 10534 11450 10590 11452
rect 10614 11450 10670 11452
rect 10374 11398 10420 11450
rect 10420 11398 10430 11450
rect 10454 11398 10484 11450
rect 10484 11398 10496 11450
rect 10496 11398 10510 11450
rect 10534 11398 10548 11450
rect 10548 11398 10560 11450
rect 10560 11398 10590 11450
rect 10614 11398 10624 11450
rect 10624 11398 10670 11450
rect 10374 11396 10430 11398
rect 10454 11396 10510 11398
rect 10534 11396 10590 11398
rect 10614 11396 10670 11398
rect 8114 2916 8170 2952
rect 9126 3576 9182 3632
rect 9402 3440 9458 3496
rect 9862 3984 9918 4040
rect 9678 3032 9734 3088
rect 8114 2896 8116 2916
rect 8116 2896 8168 2916
rect 8168 2896 8170 2916
rect 7683 2746 7739 2748
rect 7763 2746 7819 2748
rect 7843 2746 7899 2748
rect 7923 2746 7979 2748
rect 7683 2694 7729 2746
rect 7729 2694 7739 2746
rect 7763 2694 7793 2746
rect 7793 2694 7805 2746
rect 7805 2694 7819 2746
rect 7843 2694 7857 2746
rect 7857 2694 7869 2746
rect 7869 2694 7899 2746
rect 7923 2694 7933 2746
rect 7933 2694 7979 2746
rect 7683 2692 7739 2694
rect 7763 2692 7819 2694
rect 7843 2692 7899 2694
rect 7923 2692 7979 2694
rect 7470 2644 7526 2680
rect 7470 2624 7472 2644
rect 7472 2624 7524 2644
rect 7524 2624 7526 2644
rect 10046 6840 10102 6896
rect 10374 10362 10430 10364
rect 10454 10362 10510 10364
rect 10534 10362 10590 10364
rect 10614 10362 10670 10364
rect 10374 10310 10420 10362
rect 10420 10310 10430 10362
rect 10454 10310 10484 10362
rect 10484 10310 10496 10362
rect 10496 10310 10510 10362
rect 10534 10310 10548 10362
rect 10548 10310 10560 10362
rect 10560 10310 10590 10362
rect 10614 10310 10624 10362
rect 10624 10310 10670 10362
rect 10374 10308 10430 10310
rect 10454 10308 10510 10310
rect 10534 10308 10590 10310
rect 10614 10308 10670 10310
rect 11518 10920 11574 10976
rect 11034 10906 11090 10908
rect 11114 10906 11170 10908
rect 11194 10906 11250 10908
rect 11274 10906 11330 10908
rect 11034 10854 11080 10906
rect 11080 10854 11090 10906
rect 11114 10854 11144 10906
rect 11144 10854 11156 10906
rect 11156 10854 11170 10906
rect 11194 10854 11208 10906
rect 11208 10854 11220 10906
rect 11220 10854 11250 10906
rect 11274 10854 11284 10906
rect 11284 10854 11330 10906
rect 11034 10852 11090 10854
rect 11114 10852 11170 10854
rect 11194 10852 11250 10854
rect 11274 10852 11330 10854
rect 10374 9274 10430 9276
rect 10454 9274 10510 9276
rect 10534 9274 10590 9276
rect 10614 9274 10670 9276
rect 10374 9222 10420 9274
rect 10420 9222 10430 9274
rect 10454 9222 10484 9274
rect 10484 9222 10496 9274
rect 10496 9222 10510 9274
rect 10534 9222 10548 9274
rect 10548 9222 10560 9274
rect 10560 9222 10590 9274
rect 10614 9222 10624 9274
rect 10624 9222 10670 9274
rect 10374 9220 10430 9222
rect 10454 9220 10510 9222
rect 10534 9220 10590 9222
rect 10614 9220 10670 9222
rect 11034 9818 11090 9820
rect 11114 9818 11170 9820
rect 11194 9818 11250 9820
rect 11274 9818 11330 9820
rect 11034 9766 11080 9818
rect 11080 9766 11090 9818
rect 11114 9766 11144 9818
rect 11144 9766 11156 9818
rect 11156 9766 11170 9818
rect 11194 9766 11208 9818
rect 11208 9766 11220 9818
rect 11220 9766 11250 9818
rect 11274 9766 11284 9818
rect 11284 9766 11330 9818
rect 11034 9764 11090 9766
rect 11114 9764 11170 9766
rect 11194 9764 11250 9766
rect 11274 9764 11330 9766
rect 11518 9560 11574 9616
rect 11034 8730 11090 8732
rect 11114 8730 11170 8732
rect 11194 8730 11250 8732
rect 11274 8730 11330 8732
rect 11034 8678 11080 8730
rect 11080 8678 11090 8730
rect 11114 8678 11144 8730
rect 11144 8678 11156 8730
rect 11156 8678 11170 8730
rect 11194 8678 11208 8730
rect 11208 8678 11220 8730
rect 11220 8678 11250 8730
rect 11274 8678 11284 8730
rect 11284 8678 11330 8730
rect 11034 8676 11090 8678
rect 11114 8676 11170 8678
rect 11194 8676 11250 8678
rect 11274 8676 11330 8678
rect 10374 8186 10430 8188
rect 10454 8186 10510 8188
rect 10534 8186 10590 8188
rect 10614 8186 10670 8188
rect 10374 8134 10420 8186
rect 10420 8134 10430 8186
rect 10454 8134 10484 8186
rect 10484 8134 10496 8186
rect 10496 8134 10510 8186
rect 10534 8134 10548 8186
rect 10548 8134 10560 8186
rect 10560 8134 10590 8186
rect 10614 8134 10624 8186
rect 10624 8134 10670 8186
rect 10374 8132 10430 8134
rect 10454 8132 10510 8134
rect 10534 8132 10590 8134
rect 10614 8132 10670 8134
rect 10374 7098 10430 7100
rect 10454 7098 10510 7100
rect 10534 7098 10590 7100
rect 10614 7098 10670 7100
rect 10374 7046 10420 7098
rect 10420 7046 10430 7098
rect 10454 7046 10484 7098
rect 10484 7046 10496 7098
rect 10496 7046 10510 7098
rect 10534 7046 10548 7098
rect 10548 7046 10560 7098
rect 10560 7046 10590 7098
rect 10614 7046 10624 7098
rect 10624 7046 10670 7098
rect 10374 7044 10430 7046
rect 10454 7044 10510 7046
rect 10534 7044 10590 7046
rect 10614 7044 10670 7046
rect 10414 6840 10470 6896
rect 11034 7642 11090 7644
rect 11114 7642 11170 7644
rect 11194 7642 11250 7644
rect 11274 7642 11330 7644
rect 11034 7590 11080 7642
rect 11080 7590 11090 7642
rect 11114 7590 11144 7642
rect 11144 7590 11156 7642
rect 11156 7590 11170 7642
rect 11194 7590 11208 7642
rect 11208 7590 11220 7642
rect 11220 7590 11250 7642
rect 11274 7590 11284 7642
rect 11284 7590 11330 7642
rect 11034 7588 11090 7590
rect 11114 7588 11170 7590
rect 11194 7588 11250 7590
rect 11274 7588 11330 7590
rect 11518 8200 11574 8256
rect 11242 6840 11298 6896
rect 11426 6568 11482 6624
rect 11034 6554 11090 6556
rect 11114 6554 11170 6556
rect 11194 6554 11250 6556
rect 11274 6554 11330 6556
rect 11034 6502 11080 6554
rect 11080 6502 11090 6554
rect 11114 6502 11144 6554
rect 11144 6502 11156 6554
rect 11156 6502 11170 6554
rect 11194 6502 11208 6554
rect 11208 6502 11220 6554
rect 11220 6502 11250 6554
rect 11274 6502 11284 6554
rect 11284 6502 11330 6554
rect 11034 6500 11090 6502
rect 11114 6500 11170 6502
rect 11194 6500 11250 6502
rect 11274 6500 11330 6502
rect 10782 6296 10838 6352
rect 10598 6160 10654 6216
rect 10782 6160 10838 6216
rect 10374 6010 10430 6012
rect 10454 6010 10510 6012
rect 10534 6010 10590 6012
rect 10614 6010 10670 6012
rect 10374 5958 10420 6010
rect 10420 5958 10430 6010
rect 10454 5958 10484 6010
rect 10484 5958 10496 6010
rect 10496 5958 10510 6010
rect 10534 5958 10548 6010
rect 10548 5958 10560 6010
rect 10560 5958 10590 6010
rect 10614 5958 10624 6010
rect 10624 5958 10670 6010
rect 10374 5956 10430 5958
rect 10454 5956 10510 5958
rect 10534 5956 10590 5958
rect 10614 5956 10670 5958
rect 10506 5752 10562 5808
rect 10230 5616 10286 5672
rect 10374 4922 10430 4924
rect 10454 4922 10510 4924
rect 10534 4922 10590 4924
rect 10614 4922 10670 4924
rect 10374 4870 10420 4922
rect 10420 4870 10430 4922
rect 10454 4870 10484 4922
rect 10484 4870 10496 4922
rect 10496 4870 10510 4922
rect 10534 4870 10548 4922
rect 10548 4870 10560 4922
rect 10560 4870 10590 4922
rect 10614 4870 10624 4922
rect 10624 4870 10670 4922
rect 10374 4868 10430 4870
rect 10454 4868 10510 4870
rect 10534 4868 10590 4870
rect 10614 4868 10670 4870
rect 10374 3834 10430 3836
rect 10454 3834 10510 3836
rect 10534 3834 10590 3836
rect 10614 3834 10670 3836
rect 10374 3782 10420 3834
rect 10420 3782 10430 3834
rect 10454 3782 10484 3834
rect 10484 3782 10496 3834
rect 10496 3782 10510 3834
rect 10534 3782 10548 3834
rect 10548 3782 10560 3834
rect 10560 3782 10590 3834
rect 10614 3782 10624 3834
rect 10624 3782 10670 3834
rect 10374 3780 10430 3782
rect 10454 3780 10510 3782
rect 10534 3780 10590 3782
rect 10614 3780 10670 3782
rect 11334 5652 11336 5672
rect 11336 5652 11388 5672
rect 11388 5652 11390 5672
rect 11334 5616 11390 5652
rect 11034 5466 11090 5468
rect 11114 5466 11170 5468
rect 11194 5466 11250 5468
rect 11274 5466 11330 5468
rect 11034 5414 11080 5466
rect 11080 5414 11090 5466
rect 11114 5414 11144 5466
rect 11144 5414 11156 5466
rect 11156 5414 11170 5466
rect 11194 5414 11208 5466
rect 11208 5414 11220 5466
rect 11220 5414 11250 5466
rect 11274 5414 11284 5466
rect 11284 5414 11330 5466
rect 11034 5412 11090 5414
rect 11114 5412 11170 5414
rect 11194 5412 11250 5414
rect 11274 5412 11330 5414
rect 11518 5480 11574 5536
rect 11034 4378 11090 4380
rect 11114 4378 11170 4380
rect 11194 4378 11250 4380
rect 11274 4378 11330 4380
rect 11034 4326 11080 4378
rect 11080 4326 11090 4378
rect 11114 4326 11144 4378
rect 11144 4326 11156 4378
rect 11156 4326 11170 4378
rect 11194 4326 11208 4378
rect 11208 4326 11220 4378
rect 11220 4326 11250 4378
rect 11274 4326 11284 4378
rect 11284 4326 11330 4378
rect 11034 4324 11090 4326
rect 11114 4324 11170 4326
rect 11194 4324 11250 4326
rect 11274 4324 11330 4326
rect 11426 4120 11482 4176
rect 11034 3290 11090 3292
rect 11114 3290 11170 3292
rect 11194 3290 11250 3292
rect 11274 3290 11330 3292
rect 11034 3238 11080 3290
rect 11080 3238 11090 3290
rect 11114 3238 11144 3290
rect 11144 3238 11156 3290
rect 11156 3238 11170 3290
rect 11194 3238 11208 3290
rect 11208 3238 11220 3290
rect 11220 3238 11250 3290
rect 11274 3238 11284 3290
rect 11284 3238 11330 3290
rect 11034 3236 11090 3238
rect 11114 3236 11170 3238
rect 11194 3236 11250 3238
rect 11274 3236 11330 3238
rect 10374 2746 10430 2748
rect 10454 2746 10510 2748
rect 10534 2746 10590 2748
rect 10614 2746 10670 2748
rect 10374 2694 10420 2746
rect 10420 2694 10430 2746
rect 10454 2694 10484 2746
rect 10484 2694 10496 2746
rect 10496 2694 10510 2746
rect 10534 2694 10548 2746
rect 10548 2694 10560 2746
rect 10560 2694 10590 2746
rect 10614 2694 10624 2746
rect 10624 2694 10670 2746
rect 10374 2692 10430 2694
rect 10454 2692 10510 2694
rect 10534 2692 10590 2694
rect 10614 2692 10670 2694
rect 11334 2760 11390 2816
rect 5652 2202 5708 2204
rect 5732 2202 5788 2204
rect 5812 2202 5868 2204
rect 5892 2202 5948 2204
rect 5652 2150 5698 2202
rect 5698 2150 5708 2202
rect 5732 2150 5762 2202
rect 5762 2150 5774 2202
rect 5774 2150 5788 2202
rect 5812 2150 5826 2202
rect 5826 2150 5838 2202
rect 5838 2150 5868 2202
rect 5892 2150 5902 2202
rect 5902 2150 5948 2202
rect 5652 2148 5708 2150
rect 5732 2148 5788 2150
rect 5812 2148 5868 2150
rect 5892 2148 5948 2150
rect 8343 2202 8399 2204
rect 8423 2202 8479 2204
rect 8503 2202 8559 2204
rect 8583 2202 8639 2204
rect 8343 2150 8389 2202
rect 8389 2150 8399 2202
rect 8423 2150 8453 2202
rect 8453 2150 8465 2202
rect 8465 2150 8479 2202
rect 8503 2150 8517 2202
rect 8517 2150 8529 2202
rect 8529 2150 8559 2202
rect 8583 2150 8593 2202
rect 8593 2150 8639 2202
rect 8343 2148 8399 2150
rect 8423 2148 8479 2150
rect 8503 2148 8559 2150
rect 8583 2148 8639 2150
rect 11034 2202 11090 2204
rect 11114 2202 11170 2204
rect 11194 2202 11250 2204
rect 11274 2202 11330 2204
rect 11034 2150 11080 2202
rect 11080 2150 11090 2202
rect 11114 2150 11144 2202
rect 11144 2150 11156 2202
rect 11156 2150 11170 2202
rect 11194 2150 11208 2202
rect 11208 2150 11220 2202
rect 11220 2150 11250 2202
rect 11274 2150 11284 2202
rect 11284 2150 11330 2202
rect 11034 2148 11090 2150
rect 11114 2148 11170 2150
rect 11194 2148 11250 2150
rect 11274 2148 11330 2150
rect 11426 1400 11482 1456
<< metal3 >>
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 11421 13698 11487 13701
rect 12253 13698 13053 13728
rect 11421 13696 13053 13698
rect 11421 13640 11426 13696
rect 11482 13640 13053 13696
rect 11421 13638 13053 13640
rect 11421 13635 11487 13638
rect 12253 13608 13053 13638
rect 2291 12544 2607 12545
rect 2291 12480 2297 12544
rect 2361 12480 2377 12544
rect 2441 12480 2457 12544
rect 2521 12480 2537 12544
rect 2601 12480 2607 12544
rect 2291 12479 2607 12480
rect 4982 12544 5298 12545
rect 4982 12480 4988 12544
rect 5052 12480 5068 12544
rect 5132 12480 5148 12544
rect 5212 12480 5228 12544
rect 5292 12480 5298 12544
rect 4982 12479 5298 12480
rect 7673 12544 7989 12545
rect 7673 12480 7679 12544
rect 7743 12480 7759 12544
rect 7823 12480 7839 12544
rect 7903 12480 7919 12544
rect 7983 12480 7989 12544
rect 7673 12479 7989 12480
rect 10364 12544 10680 12545
rect 10364 12480 10370 12544
rect 10434 12480 10450 12544
rect 10514 12480 10530 12544
rect 10594 12480 10610 12544
rect 10674 12480 10680 12544
rect 10364 12479 10680 12480
rect 0 12338 800 12368
rect 1025 12338 1091 12341
rect 0 12336 1091 12338
rect 0 12280 1030 12336
rect 1086 12280 1091 12336
rect 0 12278 1091 12280
rect 0 12248 800 12278
rect 1025 12275 1091 12278
rect 11513 12338 11579 12341
rect 12253 12338 13053 12368
rect 11513 12336 13053 12338
rect 11513 12280 11518 12336
rect 11574 12280 13053 12336
rect 11513 12278 13053 12280
rect 11513 12275 11579 12278
rect 12253 12248 13053 12278
rect 2951 12000 3267 12001
rect 2951 11936 2957 12000
rect 3021 11936 3037 12000
rect 3101 11936 3117 12000
rect 3181 11936 3197 12000
rect 3261 11936 3267 12000
rect 2951 11935 3267 11936
rect 5642 12000 5958 12001
rect 5642 11936 5648 12000
rect 5712 11936 5728 12000
rect 5792 11936 5808 12000
rect 5872 11936 5888 12000
rect 5952 11936 5958 12000
rect 5642 11935 5958 11936
rect 8333 12000 8649 12001
rect 8333 11936 8339 12000
rect 8403 11936 8419 12000
rect 8483 11936 8499 12000
rect 8563 11936 8579 12000
rect 8643 11936 8649 12000
rect 8333 11935 8649 11936
rect 11024 12000 11340 12001
rect 11024 11936 11030 12000
rect 11094 11936 11110 12000
rect 11174 11936 11190 12000
rect 11254 11936 11270 12000
rect 11334 11936 11340 12000
rect 11024 11935 11340 11936
rect 1853 11658 1919 11661
rect 6453 11658 6519 11661
rect 1853 11656 6519 11658
rect 1853 11600 1858 11656
rect 1914 11600 6458 11656
rect 6514 11600 6519 11656
rect 1853 11598 6519 11600
rect 1853 11595 1919 11598
rect 6453 11595 6519 11598
rect 2291 11456 2607 11457
rect 2291 11392 2297 11456
rect 2361 11392 2377 11456
rect 2441 11392 2457 11456
rect 2521 11392 2537 11456
rect 2601 11392 2607 11456
rect 2291 11391 2607 11392
rect 4982 11456 5298 11457
rect 4982 11392 4988 11456
rect 5052 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5298 11456
rect 4982 11391 5298 11392
rect 7673 11456 7989 11457
rect 7673 11392 7679 11456
rect 7743 11392 7759 11456
rect 7823 11392 7839 11456
rect 7903 11392 7919 11456
rect 7983 11392 7989 11456
rect 7673 11391 7989 11392
rect 10364 11456 10680 11457
rect 10364 11392 10370 11456
rect 10434 11392 10450 11456
rect 10514 11392 10530 11456
rect 10594 11392 10610 11456
rect 10674 11392 10680 11456
rect 10364 11391 10680 11392
rect 4245 11114 4311 11117
rect 8937 11114 9003 11117
rect 4245 11112 9003 11114
rect 4245 11056 4250 11112
rect 4306 11056 8942 11112
rect 8998 11056 9003 11112
rect 4245 11054 9003 11056
rect 4245 11051 4311 11054
rect 8937 11051 9003 11054
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 11513 10978 11579 10981
rect 12253 10978 13053 11008
rect 11513 10976 13053 10978
rect 11513 10920 11518 10976
rect 11574 10920 13053 10976
rect 11513 10918 13053 10920
rect 11513 10915 11579 10918
rect 2951 10912 3267 10913
rect 2951 10848 2957 10912
rect 3021 10848 3037 10912
rect 3101 10848 3117 10912
rect 3181 10848 3197 10912
rect 3261 10848 3267 10912
rect 2951 10847 3267 10848
rect 5642 10912 5958 10913
rect 5642 10848 5648 10912
rect 5712 10848 5728 10912
rect 5792 10848 5808 10912
rect 5872 10848 5888 10912
rect 5952 10848 5958 10912
rect 5642 10847 5958 10848
rect 8333 10912 8649 10913
rect 8333 10848 8339 10912
rect 8403 10848 8419 10912
rect 8483 10848 8499 10912
rect 8563 10848 8579 10912
rect 8643 10848 8649 10912
rect 8333 10847 8649 10848
rect 11024 10912 11340 10913
rect 11024 10848 11030 10912
rect 11094 10848 11110 10912
rect 11174 10848 11190 10912
rect 11254 10848 11270 10912
rect 11334 10848 11340 10912
rect 12253 10888 13053 10918
rect 11024 10847 11340 10848
rect 2291 10368 2607 10369
rect 2291 10304 2297 10368
rect 2361 10304 2377 10368
rect 2441 10304 2457 10368
rect 2521 10304 2537 10368
rect 2601 10304 2607 10368
rect 2291 10303 2607 10304
rect 4982 10368 5298 10369
rect 4982 10304 4988 10368
rect 5052 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5298 10368
rect 4982 10303 5298 10304
rect 7673 10368 7989 10369
rect 7673 10304 7679 10368
rect 7743 10304 7759 10368
rect 7823 10304 7839 10368
rect 7903 10304 7919 10368
rect 7983 10304 7989 10368
rect 7673 10303 7989 10304
rect 10364 10368 10680 10369
rect 10364 10304 10370 10368
rect 10434 10304 10450 10368
rect 10514 10304 10530 10368
rect 10594 10304 10610 10368
rect 10674 10304 10680 10368
rect 10364 10303 10680 10304
rect 7465 9892 7531 9893
rect 7414 9828 7420 9892
rect 7484 9890 7531 9892
rect 7484 9888 7576 9890
rect 7526 9832 7576 9888
rect 7484 9830 7576 9832
rect 7484 9828 7531 9830
rect 7465 9827 7531 9828
rect 2951 9824 3267 9825
rect 2951 9760 2957 9824
rect 3021 9760 3037 9824
rect 3101 9760 3117 9824
rect 3181 9760 3197 9824
rect 3261 9760 3267 9824
rect 2951 9759 3267 9760
rect 5642 9824 5958 9825
rect 5642 9760 5648 9824
rect 5712 9760 5728 9824
rect 5792 9760 5808 9824
rect 5872 9760 5888 9824
rect 5952 9760 5958 9824
rect 5642 9759 5958 9760
rect 8333 9824 8649 9825
rect 8333 9760 8339 9824
rect 8403 9760 8419 9824
rect 8483 9760 8499 9824
rect 8563 9760 8579 9824
rect 8643 9760 8649 9824
rect 8333 9759 8649 9760
rect 11024 9824 11340 9825
rect 11024 9760 11030 9824
rect 11094 9760 11110 9824
rect 11174 9760 11190 9824
rect 11254 9760 11270 9824
rect 11334 9760 11340 9824
rect 11024 9759 11340 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 11513 9618 11579 9621
rect 12253 9618 13053 9648
rect 11513 9616 13053 9618
rect 11513 9560 11518 9616
rect 11574 9560 13053 9616
rect 11513 9558 13053 9560
rect 11513 9555 11579 9558
rect 12253 9528 13053 9558
rect 2291 9280 2607 9281
rect 2291 9216 2297 9280
rect 2361 9216 2377 9280
rect 2441 9216 2457 9280
rect 2521 9216 2537 9280
rect 2601 9216 2607 9280
rect 2291 9215 2607 9216
rect 4982 9280 5298 9281
rect 4982 9216 4988 9280
rect 5052 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5298 9280
rect 4982 9215 5298 9216
rect 7673 9280 7989 9281
rect 7673 9216 7679 9280
rect 7743 9216 7759 9280
rect 7823 9216 7839 9280
rect 7903 9216 7919 9280
rect 7983 9216 7989 9280
rect 7673 9215 7989 9216
rect 10364 9280 10680 9281
rect 10364 9216 10370 9280
rect 10434 9216 10450 9280
rect 10514 9216 10530 9280
rect 10594 9216 10610 9280
rect 10674 9216 10680 9280
rect 10364 9215 10680 9216
rect 6361 8938 6427 8941
rect 6361 8936 6562 8938
rect 6361 8880 6366 8936
rect 6422 8880 6562 8936
rect 6361 8878 6562 8880
rect 6361 8875 6427 8878
rect 2951 8736 3267 8737
rect 2951 8672 2957 8736
rect 3021 8672 3037 8736
rect 3101 8672 3117 8736
rect 3181 8672 3197 8736
rect 3261 8672 3267 8736
rect 2951 8671 3267 8672
rect 5642 8736 5958 8737
rect 5642 8672 5648 8736
rect 5712 8672 5728 8736
rect 5792 8672 5808 8736
rect 5872 8672 5888 8736
rect 5952 8672 5958 8736
rect 5642 8671 5958 8672
rect 5165 8394 5231 8397
rect 4662 8392 5231 8394
rect 4662 8336 5170 8392
rect 5226 8336 5231 8392
rect 4662 8334 5231 8336
rect 6502 8394 6562 8878
rect 8333 8736 8649 8737
rect 8333 8672 8339 8736
rect 8403 8672 8419 8736
rect 8483 8672 8499 8736
rect 8563 8672 8579 8736
rect 8643 8672 8649 8736
rect 8333 8671 8649 8672
rect 11024 8736 11340 8737
rect 11024 8672 11030 8736
rect 11094 8672 11110 8736
rect 11174 8672 11190 8736
rect 11254 8672 11270 8736
rect 11334 8672 11340 8736
rect 11024 8671 11340 8672
rect 6729 8394 6795 8397
rect 6502 8392 6795 8394
rect 6502 8336 6734 8392
rect 6790 8336 6795 8392
rect 6502 8334 6795 8336
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 2291 8192 2607 8193
rect 2291 8128 2297 8192
rect 2361 8128 2377 8192
rect 2441 8128 2457 8192
rect 2521 8128 2537 8192
rect 2601 8128 2607 8192
rect 2291 8127 2607 8128
rect 4662 7989 4722 8334
rect 5165 8331 5231 8334
rect 6729 8331 6795 8334
rect 8937 8258 9003 8261
rect 9397 8258 9463 8261
rect 8937 8256 9463 8258
rect 8937 8200 8942 8256
rect 8998 8200 9402 8256
rect 9458 8200 9463 8256
rect 8937 8198 9463 8200
rect 8937 8195 9003 8198
rect 9397 8195 9463 8198
rect 11513 8258 11579 8261
rect 12253 8258 13053 8288
rect 11513 8256 13053 8258
rect 11513 8200 11518 8256
rect 11574 8200 13053 8256
rect 11513 8198 13053 8200
rect 11513 8195 11579 8198
rect 4982 8192 5298 8193
rect 4982 8128 4988 8192
rect 5052 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5298 8192
rect 4982 8127 5298 8128
rect 7673 8192 7989 8193
rect 7673 8128 7679 8192
rect 7743 8128 7759 8192
rect 7823 8128 7839 8192
rect 7903 8128 7919 8192
rect 7983 8128 7989 8192
rect 7673 8127 7989 8128
rect 10364 8192 10680 8193
rect 10364 8128 10370 8192
rect 10434 8128 10450 8192
rect 10514 8128 10530 8192
rect 10594 8128 10610 8192
rect 10674 8128 10680 8192
rect 12253 8168 13053 8198
rect 10364 8127 10680 8128
rect 3233 7986 3299 7989
rect 3233 7984 3572 7986
rect 3233 7928 3238 7984
rect 3294 7928 3572 7984
rect 3233 7926 3572 7928
rect 3233 7923 3299 7926
rect 3512 7853 3572 7926
rect 4613 7984 4722 7989
rect 4613 7928 4618 7984
rect 4674 7928 4722 7984
rect 4613 7926 4722 7928
rect 4613 7923 4679 7926
rect 3509 7848 3575 7853
rect 3509 7792 3514 7848
rect 3570 7792 3575 7848
rect 3509 7787 3575 7792
rect 2951 7648 3267 7649
rect 2951 7584 2957 7648
rect 3021 7584 3037 7648
rect 3101 7584 3117 7648
rect 3181 7584 3197 7648
rect 3261 7584 3267 7648
rect 2951 7583 3267 7584
rect 5642 7648 5958 7649
rect 5642 7584 5648 7648
rect 5712 7584 5728 7648
rect 5792 7584 5808 7648
rect 5872 7584 5888 7648
rect 5952 7584 5958 7648
rect 5642 7583 5958 7584
rect 8333 7648 8649 7649
rect 8333 7584 8339 7648
rect 8403 7584 8419 7648
rect 8483 7584 8499 7648
rect 8563 7584 8579 7648
rect 8643 7584 8649 7648
rect 8333 7583 8649 7584
rect 11024 7648 11340 7649
rect 11024 7584 11030 7648
rect 11094 7584 11110 7648
rect 11174 7584 11190 7648
rect 11254 7584 11270 7648
rect 11334 7584 11340 7648
rect 11024 7583 11340 7584
rect 2291 7104 2607 7105
rect 2291 7040 2297 7104
rect 2361 7040 2377 7104
rect 2441 7040 2457 7104
rect 2521 7040 2537 7104
rect 2601 7040 2607 7104
rect 2291 7039 2607 7040
rect 4982 7104 5298 7105
rect 4982 7040 4988 7104
rect 5052 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5298 7104
rect 4982 7039 5298 7040
rect 7673 7104 7989 7105
rect 7673 7040 7679 7104
rect 7743 7040 7759 7104
rect 7823 7040 7839 7104
rect 7903 7040 7919 7104
rect 7983 7040 7989 7104
rect 7673 7039 7989 7040
rect 10364 7104 10680 7105
rect 10364 7040 10370 7104
rect 10434 7040 10450 7104
rect 10514 7040 10530 7104
rect 10594 7040 10610 7104
rect 10674 7040 10680 7104
rect 10364 7039 10680 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 10041 6898 10107 6901
rect 10409 6898 10475 6901
rect 10041 6896 10475 6898
rect 10041 6840 10046 6896
rect 10102 6840 10414 6896
rect 10470 6840 10475 6896
rect 10041 6838 10475 6840
rect 10041 6835 10107 6838
rect 10409 6835 10475 6838
rect 11237 6898 11303 6901
rect 12253 6898 13053 6928
rect 11237 6896 13053 6898
rect 11237 6840 11242 6896
rect 11298 6840 13053 6896
rect 11237 6838 13053 6840
rect 11237 6835 11303 6838
rect 10412 6762 10472 6835
rect 12253 6808 13053 6838
rect 10412 6702 11484 6762
rect 11424 6629 11484 6702
rect 11421 6624 11487 6629
rect 11421 6568 11426 6624
rect 11482 6568 11487 6624
rect 11421 6563 11487 6568
rect 2951 6560 3267 6561
rect 2951 6496 2957 6560
rect 3021 6496 3037 6560
rect 3101 6496 3117 6560
rect 3181 6496 3197 6560
rect 3261 6496 3267 6560
rect 2951 6495 3267 6496
rect 5642 6560 5958 6561
rect 5642 6496 5648 6560
rect 5712 6496 5728 6560
rect 5792 6496 5808 6560
rect 5872 6496 5888 6560
rect 5952 6496 5958 6560
rect 5642 6495 5958 6496
rect 8333 6560 8649 6561
rect 8333 6496 8339 6560
rect 8403 6496 8419 6560
rect 8483 6496 8499 6560
rect 8563 6496 8579 6560
rect 8643 6496 8649 6560
rect 8333 6495 8649 6496
rect 11024 6560 11340 6561
rect 11024 6496 11030 6560
rect 11094 6496 11110 6560
rect 11174 6496 11190 6560
rect 11254 6496 11270 6560
rect 11334 6496 11340 6560
rect 11024 6495 11340 6496
rect 7097 6354 7163 6357
rect 8293 6354 8359 6357
rect 7097 6352 8359 6354
rect 7097 6296 7102 6352
rect 7158 6296 8298 6352
rect 8354 6296 8359 6352
rect 7097 6294 8359 6296
rect 7097 6291 7163 6294
rect 8293 6291 8359 6294
rect 10777 6354 10843 6357
rect 10777 6352 10978 6354
rect 10777 6296 10782 6352
rect 10838 6296 10978 6352
rect 10777 6294 10978 6296
rect 10777 6291 10843 6294
rect 3601 6218 3667 6221
rect 7649 6218 7715 6221
rect 3601 6216 7715 6218
rect 3601 6160 3606 6216
rect 3662 6160 7654 6216
rect 7710 6160 7715 6216
rect 3601 6158 7715 6160
rect 3601 6155 3667 6158
rect 7649 6155 7715 6158
rect 10593 6218 10659 6221
rect 10777 6218 10843 6221
rect 10593 6216 10843 6218
rect 10593 6160 10598 6216
rect 10654 6160 10782 6216
rect 10838 6160 10843 6216
rect 10593 6158 10843 6160
rect 10593 6155 10659 6158
rect 10777 6155 10843 6158
rect 5625 6082 5691 6085
rect 6729 6082 6795 6085
rect 5625 6080 6795 6082
rect 5625 6024 5630 6080
rect 5686 6024 6734 6080
rect 6790 6024 6795 6080
rect 5625 6022 6795 6024
rect 5625 6019 5691 6022
rect 6729 6019 6795 6022
rect 2291 6016 2607 6017
rect 2291 5952 2297 6016
rect 2361 5952 2377 6016
rect 2441 5952 2457 6016
rect 2521 5952 2537 6016
rect 2601 5952 2607 6016
rect 2291 5951 2607 5952
rect 4982 6016 5298 6017
rect 4982 5952 4988 6016
rect 5052 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5298 6016
rect 4982 5951 5298 5952
rect 7673 6016 7989 6017
rect 7673 5952 7679 6016
rect 7743 5952 7759 6016
rect 7823 5952 7839 6016
rect 7903 5952 7919 6016
rect 7983 5952 7989 6016
rect 7673 5951 7989 5952
rect 10364 6016 10680 6017
rect 10364 5952 10370 6016
rect 10434 5952 10450 6016
rect 10514 5952 10530 6016
rect 10594 5952 10610 6016
rect 10674 5952 10680 6016
rect 10364 5951 10680 5952
rect 10501 5810 10567 5813
rect 10918 5810 10978 6294
rect 10501 5808 10978 5810
rect 10501 5752 10506 5808
rect 10562 5752 10978 5808
rect 10501 5750 10978 5752
rect 10501 5747 10567 5750
rect 10225 5674 10291 5677
rect 11329 5674 11395 5677
rect 10225 5672 11395 5674
rect 10225 5616 10230 5672
rect 10286 5616 11334 5672
rect 11390 5616 11395 5672
rect 10225 5614 11395 5616
rect 10225 5611 10291 5614
rect 11329 5611 11395 5614
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 11513 5538 11579 5541
rect 12253 5538 13053 5568
rect 11513 5536 13053 5538
rect 11513 5480 11518 5536
rect 11574 5480 13053 5536
rect 11513 5478 13053 5480
rect 11513 5475 11579 5478
rect 2951 5472 3267 5473
rect 2951 5408 2957 5472
rect 3021 5408 3037 5472
rect 3101 5408 3117 5472
rect 3181 5408 3197 5472
rect 3261 5408 3267 5472
rect 2951 5407 3267 5408
rect 5642 5472 5958 5473
rect 5642 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5958 5472
rect 5642 5407 5958 5408
rect 8333 5472 8649 5473
rect 8333 5408 8339 5472
rect 8403 5408 8419 5472
rect 8483 5408 8499 5472
rect 8563 5408 8579 5472
rect 8643 5408 8649 5472
rect 8333 5407 8649 5408
rect 11024 5472 11340 5473
rect 11024 5408 11030 5472
rect 11094 5408 11110 5472
rect 11174 5408 11190 5472
rect 11254 5408 11270 5472
rect 11334 5408 11340 5472
rect 12253 5448 13053 5478
rect 11024 5407 11340 5408
rect 1669 5266 1735 5269
rect 5441 5266 5507 5269
rect 6361 5266 6427 5269
rect 1669 5264 6427 5266
rect 1669 5208 1674 5264
rect 1730 5208 5446 5264
rect 5502 5208 6366 5264
rect 6422 5208 6427 5264
rect 1669 5206 6427 5208
rect 1669 5203 1735 5206
rect 5441 5203 5507 5206
rect 6361 5203 6427 5206
rect 7281 5266 7347 5269
rect 8569 5266 8635 5269
rect 7281 5264 8635 5266
rect 7281 5208 7286 5264
rect 7342 5208 8574 5264
rect 8630 5208 8635 5264
rect 7281 5206 8635 5208
rect 7281 5203 7347 5206
rect 8569 5203 8635 5206
rect 2291 4928 2607 4929
rect 2291 4864 2297 4928
rect 2361 4864 2377 4928
rect 2441 4864 2457 4928
rect 2521 4864 2537 4928
rect 2601 4864 2607 4928
rect 2291 4863 2607 4864
rect 4982 4928 5298 4929
rect 4982 4864 4988 4928
rect 5052 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5298 4928
rect 4982 4863 5298 4864
rect 7673 4928 7989 4929
rect 7673 4864 7679 4928
rect 7743 4864 7759 4928
rect 7823 4864 7839 4928
rect 7903 4864 7919 4928
rect 7983 4864 7989 4928
rect 7673 4863 7989 4864
rect 10364 4928 10680 4929
rect 10364 4864 10370 4928
rect 10434 4864 10450 4928
rect 10514 4864 10530 4928
rect 10594 4864 10610 4928
rect 10674 4864 10680 4928
rect 10364 4863 10680 4864
rect 5809 4722 5875 4725
rect 6913 4722 6979 4725
rect 5809 4720 6979 4722
rect 5809 4664 5814 4720
rect 5870 4664 6918 4720
rect 6974 4664 6979 4720
rect 5809 4662 6979 4664
rect 5809 4659 5875 4662
rect 6913 4659 6979 4662
rect 7833 4722 7899 4725
rect 8017 4722 8083 4725
rect 7833 4720 8083 4722
rect 7833 4664 7838 4720
rect 7894 4664 8022 4720
rect 8078 4664 8083 4720
rect 7833 4662 8083 4664
rect 7833 4659 7899 4662
rect 8017 4659 8083 4662
rect 3325 4586 3391 4589
rect 6177 4586 6243 4589
rect 3325 4584 6243 4586
rect 3325 4528 3330 4584
rect 3386 4528 6182 4584
rect 6238 4528 6243 4584
rect 3325 4526 6243 4528
rect 3325 4523 3391 4526
rect 6177 4523 6243 4526
rect 2951 4384 3267 4385
rect 2951 4320 2957 4384
rect 3021 4320 3037 4384
rect 3101 4320 3117 4384
rect 3181 4320 3197 4384
rect 3261 4320 3267 4384
rect 2951 4319 3267 4320
rect 5642 4384 5958 4385
rect 5642 4320 5648 4384
rect 5712 4320 5728 4384
rect 5792 4320 5808 4384
rect 5872 4320 5888 4384
rect 5952 4320 5958 4384
rect 5642 4319 5958 4320
rect 8333 4384 8649 4385
rect 8333 4320 8339 4384
rect 8403 4320 8419 4384
rect 8483 4320 8499 4384
rect 8563 4320 8579 4384
rect 8643 4320 8649 4384
rect 8333 4319 8649 4320
rect 11024 4384 11340 4385
rect 11024 4320 11030 4384
rect 11094 4320 11110 4384
rect 11174 4320 11190 4384
rect 11254 4320 11270 4384
rect 11334 4320 11340 4384
rect 11024 4319 11340 4320
rect 0 4178 800 4208
rect 1301 4178 1367 4181
rect 0 4176 1367 4178
rect 0 4120 1306 4176
rect 1362 4120 1367 4176
rect 0 4118 1367 4120
rect 0 4088 800 4118
rect 1301 4115 1367 4118
rect 11421 4178 11487 4181
rect 12253 4178 13053 4208
rect 11421 4176 13053 4178
rect 11421 4120 11426 4176
rect 11482 4120 13053 4176
rect 11421 4118 13053 4120
rect 11421 4115 11487 4118
rect 12253 4088 13053 4118
rect 1577 4042 1643 4045
rect 6269 4042 6335 4045
rect 9857 4042 9923 4045
rect 1577 4040 6335 4042
rect 1577 3984 1582 4040
rect 1638 3984 6274 4040
rect 6330 3984 6335 4040
rect 1577 3982 6335 3984
rect 1577 3979 1643 3982
rect 6269 3979 6335 3982
rect 7054 4040 9923 4042
rect 7054 3984 9862 4040
rect 9918 3984 9923 4040
rect 7054 3982 9923 3984
rect 6177 3906 6243 3909
rect 7054 3906 7114 3982
rect 9857 3979 9923 3982
rect 6177 3904 7114 3906
rect 6177 3848 6182 3904
rect 6238 3848 7114 3904
rect 6177 3846 7114 3848
rect 6177 3843 6243 3846
rect 2291 3840 2607 3841
rect 2291 3776 2297 3840
rect 2361 3776 2377 3840
rect 2441 3776 2457 3840
rect 2521 3776 2537 3840
rect 2601 3776 2607 3840
rect 2291 3775 2607 3776
rect 4982 3840 5298 3841
rect 4982 3776 4988 3840
rect 5052 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5298 3840
rect 4982 3775 5298 3776
rect 7673 3840 7989 3841
rect 7673 3776 7679 3840
rect 7743 3776 7759 3840
rect 7823 3776 7839 3840
rect 7903 3776 7919 3840
rect 7983 3776 7989 3840
rect 7673 3775 7989 3776
rect 10364 3840 10680 3841
rect 10364 3776 10370 3840
rect 10434 3776 10450 3840
rect 10514 3776 10530 3840
rect 10594 3776 10610 3840
rect 10674 3776 10680 3840
rect 10364 3775 10680 3776
rect 6729 3634 6795 3637
rect 7097 3634 7163 3637
rect 9121 3634 9187 3637
rect 6729 3632 9187 3634
rect 6729 3576 6734 3632
rect 6790 3576 7102 3632
rect 7158 3576 9126 3632
rect 9182 3576 9187 3632
rect 6729 3574 9187 3576
rect 6729 3571 6795 3574
rect 7097 3571 7163 3574
rect 9121 3571 9187 3574
rect 4245 3498 4311 3501
rect 6821 3498 6887 3501
rect 9397 3498 9463 3501
rect 4245 3496 9463 3498
rect 4245 3440 4250 3496
rect 4306 3440 6826 3496
rect 6882 3440 9402 3496
rect 9458 3440 9463 3496
rect 4245 3438 9463 3440
rect 4245 3435 4311 3438
rect 6821 3435 6887 3438
rect 9397 3435 9463 3438
rect 6453 3362 6519 3365
rect 7373 3362 7439 3365
rect 6453 3360 7439 3362
rect 6453 3304 6458 3360
rect 6514 3304 7378 3360
rect 7434 3304 7439 3360
rect 6453 3302 7439 3304
rect 6453 3299 6519 3302
rect 7373 3299 7439 3302
rect 2951 3296 3267 3297
rect 2951 3232 2957 3296
rect 3021 3232 3037 3296
rect 3101 3232 3117 3296
rect 3181 3232 3197 3296
rect 3261 3232 3267 3296
rect 2951 3231 3267 3232
rect 5642 3296 5958 3297
rect 5642 3232 5648 3296
rect 5712 3232 5728 3296
rect 5792 3232 5808 3296
rect 5872 3232 5888 3296
rect 5952 3232 5958 3296
rect 5642 3231 5958 3232
rect 8333 3296 8649 3297
rect 8333 3232 8339 3296
rect 8403 3232 8419 3296
rect 8483 3232 8499 3296
rect 8563 3232 8579 3296
rect 8643 3232 8649 3296
rect 8333 3231 8649 3232
rect 11024 3296 11340 3297
rect 11024 3232 11030 3296
rect 11094 3232 11110 3296
rect 11174 3232 11190 3296
rect 11254 3232 11270 3296
rect 11334 3232 11340 3296
rect 11024 3231 11340 3232
rect 2589 3090 2655 3093
rect 5809 3090 5875 3093
rect 9673 3090 9739 3093
rect 2589 3088 9739 3090
rect 2589 3032 2594 3088
rect 2650 3032 5814 3088
rect 5870 3032 9678 3088
rect 9734 3032 9739 3088
rect 2589 3030 9739 3032
rect 2589 3027 2655 3030
rect 5809 3027 5875 3030
rect 9673 3027 9739 3030
rect 2313 2954 2379 2957
rect 5901 2954 5967 2957
rect 2313 2952 5967 2954
rect 2313 2896 2318 2952
rect 2374 2896 5906 2952
rect 5962 2896 5967 2952
rect 2313 2894 5967 2896
rect 2313 2891 2379 2894
rect 5901 2891 5967 2894
rect 6361 2954 6427 2957
rect 8109 2954 8175 2957
rect 6361 2952 8175 2954
rect 6361 2896 6366 2952
rect 6422 2896 8114 2952
rect 8170 2896 8175 2952
rect 6361 2894 8175 2896
rect 6361 2891 6427 2894
rect 8109 2891 8175 2894
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 11329 2818 11395 2821
rect 12253 2818 13053 2848
rect 11329 2816 13053 2818
rect 11329 2760 11334 2816
rect 11390 2760 13053 2816
rect 11329 2758 13053 2760
rect 11329 2755 11395 2758
rect 2291 2752 2607 2753
rect 2291 2688 2297 2752
rect 2361 2688 2377 2752
rect 2441 2688 2457 2752
rect 2521 2688 2537 2752
rect 2601 2688 2607 2752
rect 2291 2687 2607 2688
rect 4982 2752 5298 2753
rect 4982 2688 4988 2752
rect 5052 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5298 2752
rect 4982 2687 5298 2688
rect 7673 2752 7989 2753
rect 7673 2688 7679 2752
rect 7743 2688 7759 2752
rect 7823 2688 7839 2752
rect 7903 2688 7919 2752
rect 7983 2688 7989 2752
rect 7673 2687 7989 2688
rect 10364 2752 10680 2753
rect 10364 2688 10370 2752
rect 10434 2688 10450 2752
rect 10514 2688 10530 2752
rect 10594 2688 10610 2752
rect 10674 2688 10680 2752
rect 12253 2728 13053 2758
rect 10364 2687 10680 2688
rect 7465 2684 7531 2685
rect 7414 2620 7420 2684
rect 7484 2682 7531 2684
rect 7484 2680 7576 2682
rect 7526 2624 7576 2680
rect 7484 2622 7576 2624
rect 7484 2620 7531 2622
rect 7465 2619 7531 2620
rect 2951 2208 3267 2209
rect 2951 2144 2957 2208
rect 3021 2144 3037 2208
rect 3101 2144 3117 2208
rect 3181 2144 3197 2208
rect 3261 2144 3267 2208
rect 2951 2143 3267 2144
rect 5642 2208 5958 2209
rect 5642 2144 5648 2208
rect 5712 2144 5728 2208
rect 5792 2144 5808 2208
rect 5872 2144 5888 2208
rect 5952 2144 5958 2208
rect 5642 2143 5958 2144
rect 8333 2208 8649 2209
rect 8333 2144 8339 2208
rect 8403 2144 8419 2208
rect 8483 2144 8499 2208
rect 8563 2144 8579 2208
rect 8643 2144 8649 2208
rect 8333 2143 8649 2144
rect 11024 2208 11340 2209
rect 11024 2144 11030 2208
rect 11094 2144 11110 2208
rect 11174 2144 11190 2208
rect 11254 2144 11270 2208
rect 11334 2144 11340 2208
rect 11024 2143 11340 2144
rect 0 1458 800 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 800 1398
rect 1393 1395 1459 1398
rect 11421 1458 11487 1461
rect 12253 1458 13053 1488
rect 11421 1456 13053 1458
rect 11421 1400 11426 1456
rect 11482 1400 13053 1456
rect 11421 1398 13053 1400
rect 11421 1395 11487 1398
rect 12253 1368 13053 1398
<< via3 >>
rect 2297 12540 2361 12544
rect 2297 12484 2301 12540
rect 2301 12484 2357 12540
rect 2357 12484 2361 12540
rect 2297 12480 2361 12484
rect 2377 12540 2441 12544
rect 2377 12484 2381 12540
rect 2381 12484 2437 12540
rect 2437 12484 2441 12540
rect 2377 12480 2441 12484
rect 2457 12540 2521 12544
rect 2457 12484 2461 12540
rect 2461 12484 2517 12540
rect 2517 12484 2521 12540
rect 2457 12480 2521 12484
rect 2537 12540 2601 12544
rect 2537 12484 2541 12540
rect 2541 12484 2597 12540
rect 2597 12484 2601 12540
rect 2537 12480 2601 12484
rect 4988 12540 5052 12544
rect 4988 12484 4992 12540
rect 4992 12484 5048 12540
rect 5048 12484 5052 12540
rect 4988 12480 5052 12484
rect 5068 12540 5132 12544
rect 5068 12484 5072 12540
rect 5072 12484 5128 12540
rect 5128 12484 5132 12540
rect 5068 12480 5132 12484
rect 5148 12540 5212 12544
rect 5148 12484 5152 12540
rect 5152 12484 5208 12540
rect 5208 12484 5212 12540
rect 5148 12480 5212 12484
rect 5228 12540 5292 12544
rect 5228 12484 5232 12540
rect 5232 12484 5288 12540
rect 5288 12484 5292 12540
rect 5228 12480 5292 12484
rect 7679 12540 7743 12544
rect 7679 12484 7683 12540
rect 7683 12484 7739 12540
rect 7739 12484 7743 12540
rect 7679 12480 7743 12484
rect 7759 12540 7823 12544
rect 7759 12484 7763 12540
rect 7763 12484 7819 12540
rect 7819 12484 7823 12540
rect 7759 12480 7823 12484
rect 7839 12540 7903 12544
rect 7839 12484 7843 12540
rect 7843 12484 7899 12540
rect 7899 12484 7903 12540
rect 7839 12480 7903 12484
rect 7919 12540 7983 12544
rect 7919 12484 7923 12540
rect 7923 12484 7979 12540
rect 7979 12484 7983 12540
rect 7919 12480 7983 12484
rect 10370 12540 10434 12544
rect 10370 12484 10374 12540
rect 10374 12484 10430 12540
rect 10430 12484 10434 12540
rect 10370 12480 10434 12484
rect 10450 12540 10514 12544
rect 10450 12484 10454 12540
rect 10454 12484 10510 12540
rect 10510 12484 10514 12540
rect 10450 12480 10514 12484
rect 10530 12540 10594 12544
rect 10530 12484 10534 12540
rect 10534 12484 10590 12540
rect 10590 12484 10594 12540
rect 10530 12480 10594 12484
rect 10610 12540 10674 12544
rect 10610 12484 10614 12540
rect 10614 12484 10670 12540
rect 10670 12484 10674 12540
rect 10610 12480 10674 12484
rect 2957 11996 3021 12000
rect 2957 11940 2961 11996
rect 2961 11940 3017 11996
rect 3017 11940 3021 11996
rect 2957 11936 3021 11940
rect 3037 11996 3101 12000
rect 3037 11940 3041 11996
rect 3041 11940 3097 11996
rect 3097 11940 3101 11996
rect 3037 11936 3101 11940
rect 3117 11996 3181 12000
rect 3117 11940 3121 11996
rect 3121 11940 3177 11996
rect 3177 11940 3181 11996
rect 3117 11936 3181 11940
rect 3197 11996 3261 12000
rect 3197 11940 3201 11996
rect 3201 11940 3257 11996
rect 3257 11940 3261 11996
rect 3197 11936 3261 11940
rect 5648 11996 5712 12000
rect 5648 11940 5652 11996
rect 5652 11940 5708 11996
rect 5708 11940 5712 11996
rect 5648 11936 5712 11940
rect 5728 11996 5792 12000
rect 5728 11940 5732 11996
rect 5732 11940 5788 11996
rect 5788 11940 5792 11996
rect 5728 11936 5792 11940
rect 5808 11996 5872 12000
rect 5808 11940 5812 11996
rect 5812 11940 5868 11996
rect 5868 11940 5872 11996
rect 5808 11936 5872 11940
rect 5888 11996 5952 12000
rect 5888 11940 5892 11996
rect 5892 11940 5948 11996
rect 5948 11940 5952 11996
rect 5888 11936 5952 11940
rect 8339 11996 8403 12000
rect 8339 11940 8343 11996
rect 8343 11940 8399 11996
rect 8399 11940 8403 11996
rect 8339 11936 8403 11940
rect 8419 11996 8483 12000
rect 8419 11940 8423 11996
rect 8423 11940 8479 11996
rect 8479 11940 8483 11996
rect 8419 11936 8483 11940
rect 8499 11996 8563 12000
rect 8499 11940 8503 11996
rect 8503 11940 8559 11996
rect 8559 11940 8563 11996
rect 8499 11936 8563 11940
rect 8579 11996 8643 12000
rect 8579 11940 8583 11996
rect 8583 11940 8639 11996
rect 8639 11940 8643 11996
rect 8579 11936 8643 11940
rect 11030 11996 11094 12000
rect 11030 11940 11034 11996
rect 11034 11940 11090 11996
rect 11090 11940 11094 11996
rect 11030 11936 11094 11940
rect 11110 11996 11174 12000
rect 11110 11940 11114 11996
rect 11114 11940 11170 11996
rect 11170 11940 11174 11996
rect 11110 11936 11174 11940
rect 11190 11996 11254 12000
rect 11190 11940 11194 11996
rect 11194 11940 11250 11996
rect 11250 11940 11254 11996
rect 11190 11936 11254 11940
rect 11270 11996 11334 12000
rect 11270 11940 11274 11996
rect 11274 11940 11330 11996
rect 11330 11940 11334 11996
rect 11270 11936 11334 11940
rect 2297 11452 2361 11456
rect 2297 11396 2301 11452
rect 2301 11396 2357 11452
rect 2357 11396 2361 11452
rect 2297 11392 2361 11396
rect 2377 11452 2441 11456
rect 2377 11396 2381 11452
rect 2381 11396 2437 11452
rect 2437 11396 2441 11452
rect 2377 11392 2441 11396
rect 2457 11452 2521 11456
rect 2457 11396 2461 11452
rect 2461 11396 2517 11452
rect 2517 11396 2521 11452
rect 2457 11392 2521 11396
rect 2537 11452 2601 11456
rect 2537 11396 2541 11452
rect 2541 11396 2597 11452
rect 2597 11396 2601 11452
rect 2537 11392 2601 11396
rect 4988 11452 5052 11456
rect 4988 11396 4992 11452
rect 4992 11396 5048 11452
rect 5048 11396 5052 11452
rect 4988 11392 5052 11396
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 7679 11452 7743 11456
rect 7679 11396 7683 11452
rect 7683 11396 7739 11452
rect 7739 11396 7743 11452
rect 7679 11392 7743 11396
rect 7759 11452 7823 11456
rect 7759 11396 7763 11452
rect 7763 11396 7819 11452
rect 7819 11396 7823 11452
rect 7759 11392 7823 11396
rect 7839 11452 7903 11456
rect 7839 11396 7843 11452
rect 7843 11396 7899 11452
rect 7899 11396 7903 11452
rect 7839 11392 7903 11396
rect 7919 11452 7983 11456
rect 7919 11396 7923 11452
rect 7923 11396 7979 11452
rect 7979 11396 7983 11452
rect 7919 11392 7983 11396
rect 10370 11452 10434 11456
rect 10370 11396 10374 11452
rect 10374 11396 10430 11452
rect 10430 11396 10434 11452
rect 10370 11392 10434 11396
rect 10450 11452 10514 11456
rect 10450 11396 10454 11452
rect 10454 11396 10510 11452
rect 10510 11396 10514 11452
rect 10450 11392 10514 11396
rect 10530 11452 10594 11456
rect 10530 11396 10534 11452
rect 10534 11396 10590 11452
rect 10590 11396 10594 11452
rect 10530 11392 10594 11396
rect 10610 11452 10674 11456
rect 10610 11396 10614 11452
rect 10614 11396 10670 11452
rect 10670 11396 10674 11452
rect 10610 11392 10674 11396
rect 2957 10908 3021 10912
rect 2957 10852 2961 10908
rect 2961 10852 3017 10908
rect 3017 10852 3021 10908
rect 2957 10848 3021 10852
rect 3037 10908 3101 10912
rect 3037 10852 3041 10908
rect 3041 10852 3097 10908
rect 3097 10852 3101 10908
rect 3037 10848 3101 10852
rect 3117 10908 3181 10912
rect 3117 10852 3121 10908
rect 3121 10852 3177 10908
rect 3177 10852 3181 10908
rect 3117 10848 3181 10852
rect 3197 10908 3261 10912
rect 3197 10852 3201 10908
rect 3201 10852 3257 10908
rect 3257 10852 3261 10908
rect 3197 10848 3261 10852
rect 5648 10908 5712 10912
rect 5648 10852 5652 10908
rect 5652 10852 5708 10908
rect 5708 10852 5712 10908
rect 5648 10848 5712 10852
rect 5728 10908 5792 10912
rect 5728 10852 5732 10908
rect 5732 10852 5788 10908
rect 5788 10852 5792 10908
rect 5728 10848 5792 10852
rect 5808 10908 5872 10912
rect 5808 10852 5812 10908
rect 5812 10852 5868 10908
rect 5868 10852 5872 10908
rect 5808 10848 5872 10852
rect 5888 10908 5952 10912
rect 5888 10852 5892 10908
rect 5892 10852 5948 10908
rect 5948 10852 5952 10908
rect 5888 10848 5952 10852
rect 8339 10908 8403 10912
rect 8339 10852 8343 10908
rect 8343 10852 8399 10908
rect 8399 10852 8403 10908
rect 8339 10848 8403 10852
rect 8419 10908 8483 10912
rect 8419 10852 8423 10908
rect 8423 10852 8479 10908
rect 8479 10852 8483 10908
rect 8419 10848 8483 10852
rect 8499 10908 8563 10912
rect 8499 10852 8503 10908
rect 8503 10852 8559 10908
rect 8559 10852 8563 10908
rect 8499 10848 8563 10852
rect 8579 10908 8643 10912
rect 8579 10852 8583 10908
rect 8583 10852 8639 10908
rect 8639 10852 8643 10908
rect 8579 10848 8643 10852
rect 11030 10908 11094 10912
rect 11030 10852 11034 10908
rect 11034 10852 11090 10908
rect 11090 10852 11094 10908
rect 11030 10848 11094 10852
rect 11110 10908 11174 10912
rect 11110 10852 11114 10908
rect 11114 10852 11170 10908
rect 11170 10852 11174 10908
rect 11110 10848 11174 10852
rect 11190 10908 11254 10912
rect 11190 10852 11194 10908
rect 11194 10852 11250 10908
rect 11250 10852 11254 10908
rect 11190 10848 11254 10852
rect 11270 10908 11334 10912
rect 11270 10852 11274 10908
rect 11274 10852 11330 10908
rect 11330 10852 11334 10908
rect 11270 10848 11334 10852
rect 2297 10364 2361 10368
rect 2297 10308 2301 10364
rect 2301 10308 2357 10364
rect 2357 10308 2361 10364
rect 2297 10304 2361 10308
rect 2377 10364 2441 10368
rect 2377 10308 2381 10364
rect 2381 10308 2437 10364
rect 2437 10308 2441 10364
rect 2377 10304 2441 10308
rect 2457 10364 2521 10368
rect 2457 10308 2461 10364
rect 2461 10308 2517 10364
rect 2517 10308 2521 10364
rect 2457 10304 2521 10308
rect 2537 10364 2601 10368
rect 2537 10308 2541 10364
rect 2541 10308 2597 10364
rect 2597 10308 2601 10364
rect 2537 10304 2601 10308
rect 4988 10364 5052 10368
rect 4988 10308 4992 10364
rect 4992 10308 5048 10364
rect 5048 10308 5052 10364
rect 4988 10304 5052 10308
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 7679 10364 7743 10368
rect 7679 10308 7683 10364
rect 7683 10308 7739 10364
rect 7739 10308 7743 10364
rect 7679 10304 7743 10308
rect 7759 10364 7823 10368
rect 7759 10308 7763 10364
rect 7763 10308 7819 10364
rect 7819 10308 7823 10364
rect 7759 10304 7823 10308
rect 7839 10364 7903 10368
rect 7839 10308 7843 10364
rect 7843 10308 7899 10364
rect 7899 10308 7903 10364
rect 7839 10304 7903 10308
rect 7919 10364 7983 10368
rect 7919 10308 7923 10364
rect 7923 10308 7979 10364
rect 7979 10308 7983 10364
rect 7919 10304 7983 10308
rect 10370 10364 10434 10368
rect 10370 10308 10374 10364
rect 10374 10308 10430 10364
rect 10430 10308 10434 10364
rect 10370 10304 10434 10308
rect 10450 10364 10514 10368
rect 10450 10308 10454 10364
rect 10454 10308 10510 10364
rect 10510 10308 10514 10364
rect 10450 10304 10514 10308
rect 10530 10364 10594 10368
rect 10530 10308 10534 10364
rect 10534 10308 10590 10364
rect 10590 10308 10594 10364
rect 10530 10304 10594 10308
rect 10610 10364 10674 10368
rect 10610 10308 10614 10364
rect 10614 10308 10670 10364
rect 10670 10308 10674 10364
rect 10610 10304 10674 10308
rect 7420 9888 7484 9892
rect 7420 9832 7470 9888
rect 7470 9832 7484 9888
rect 7420 9828 7484 9832
rect 2957 9820 3021 9824
rect 2957 9764 2961 9820
rect 2961 9764 3017 9820
rect 3017 9764 3021 9820
rect 2957 9760 3021 9764
rect 3037 9820 3101 9824
rect 3037 9764 3041 9820
rect 3041 9764 3097 9820
rect 3097 9764 3101 9820
rect 3037 9760 3101 9764
rect 3117 9820 3181 9824
rect 3117 9764 3121 9820
rect 3121 9764 3177 9820
rect 3177 9764 3181 9820
rect 3117 9760 3181 9764
rect 3197 9820 3261 9824
rect 3197 9764 3201 9820
rect 3201 9764 3257 9820
rect 3257 9764 3261 9820
rect 3197 9760 3261 9764
rect 5648 9820 5712 9824
rect 5648 9764 5652 9820
rect 5652 9764 5708 9820
rect 5708 9764 5712 9820
rect 5648 9760 5712 9764
rect 5728 9820 5792 9824
rect 5728 9764 5732 9820
rect 5732 9764 5788 9820
rect 5788 9764 5792 9820
rect 5728 9760 5792 9764
rect 5808 9820 5872 9824
rect 5808 9764 5812 9820
rect 5812 9764 5868 9820
rect 5868 9764 5872 9820
rect 5808 9760 5872 9764
rect 5888 9820 5952 9824
rect 5888 9764 5892 9820
rect 5892 9764 5948 9820
rect 5948 9764 5952 9820
rect 5888 9760 5952 9764
rect 8339 9820 8403 9824
rect 8339 9764 8343 9820
rect 8343 9764 8399 9820
rect 8399 9764 8403 9820
rect 8339 9760 8403 9764
rect 8419 9820 8483 9824
rect 8419 9764 8423 9820
rect 8423 9764 8479 9820
rect 8479 9764 8483 9820
rect 8419 9760 8483 9764
rect 8499 9820 8563 9824
rect 8499 9764 8503 9820
rect 8503 9764 8559 9820
rect 8559 9764 8563 9820
rect 8499 9760 8563 9764
rect 8579 9820 8643 9824
rect 8579 9764 8583 9820
rect 8583 9764 8639 9820
rect 8639 9764 8643 9820
rect 8579 9760 8643 9764
rect 11030 9820 11094 9824
rect 11030 9764 11034 9820
rect 11034 9764 11090 9820
rect 11090 9764 11094 9820
rect 11030 9760 11094 9764
rect 11110 9820 11174 9824
rect 11110 9764 11114 9820
rect 11114 9764 11170 9820
rect 11170 9764 11174 9820
rect 11110 9760 11174 9764
rect 11190 9820 11254 9824
rect 11190 9764 11194 9820
rect 11194 9764 11250 9820
rect 11250 9764 11254 9820
rect 11190 9760 11254 9764
rect 11270 9820 11334 9824
rect 11270 9764 11274 9820
rect 11274 9764 11330 9820
rect 11330 9764 11334 9820
rect 11270 9760 11334 9764
rect 2297 9276 2361 9280
rect 2297 9220 2301 9276
rect 2301 9220 2357 9276
rect 2357 9220 2361 9276
rect 2297 9216 2361 9220
rect 2377 9276 2441 9280
rect 2377 9220 2381 9276
rect 2381 9220 2437 9276
rect 2437 9220 2441 9276
rect 2377 9216 2441 9220
rect 2457 9276 2521 9280
rect 2457 9220 2461 9276
rect 2461 9220 2517 9276
rect 2517 9220 2521 9276
rect 2457 9216 2521 9220
rect 2537 9276 2601 9280
rect 2537 9220 2541 9276
rect 2541 9220 2597 9276
rect 2597 9220 2601 9276
rect 2537 9216 2601 9220
rect 4988 9276 5052 9280
rect 4988 9220 4992 9276
rect 4992 9220 5048 9276
rect 5048 9220 5052 9276
rect 4988 9216 5052 9220
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 7679 9276 7743 9280
rect 7679 9220 7683 9276
rect 7683 9220 7739 9276
rect 7739 9220 7743 9276
rect 7679 9216 7743 9220
rect 7759 9276 7823 9280
rect 7759 9220 7763 9276
rect 7763 9220 7819 9276
rect 7819 9220 7823 9276
rect 7759 9216 7823 9220
rect 7839 9276 7903 9280
rect 7839 9220 7843 9276
rect 7843 9220 7899 9276
rect 7899 9220 7903 9276
rect 7839 9216 7903 9220
rect 7919 9276 7983 9280
rect 7919 9220 7923 9276
rect 7923 9220 7979 9276
rect 7979 9220 7983 9276
rect 7919 9216 7983 9220
rect 10370 9276 10434 9280
rect 10370 9220 10374 9276
rect 10374 9220 10430 9276
rect 10430 9220 10434 9276
rect 10370 9216 10434 9220
rect 10450 9276 10514 9280
rect 10450 9220 10454 9276
rect 10454 9220 10510 9276
rect 10510 9220 10514 9276
rect 10450 9216 10514 9220
rect 10530 9276 10594 9280
rect 10530 9220 10534 9276
rect 10534 9220 10590 9276
rect 10590 9220 10594 9276
rect 10530 9216 10594 9220
rect 10610 9276 10674 9280
rect 10610 9220 10614 9276
rect 10614 9220 10670 9276
rect 10670 9220 10674 9276
rect 10610 9216 10674 9220
rect 2957 8732 3021 8736
rect 2957 8676 2961 8732
rect 2961 8676 3017 8732
rect 3017 8676 3021 8732
rect 2957 8672 3021 8676
rect 3037 8732 3101 8736
rect 3037 8676 3041 8732
rect 3041 8676 3097 8732
rect 3097 8676 3101 8732
rect 3037 8672 3101 8676
rect 3117 8732 3181 8736
rect 3117 8676 3121 8732
rect 3121 8676 3177 8732
rect 3177 8676 3181 8732
rect 3117 8672 3181 8676
rect 3197 8732 3261 8736
rect 3197 8676 3201 8732
rect 3201 8676 3257 8732
rect 3257 8676 3261 8732
rect 3197 8672 3261 8676
rect 5648 8732 5712 8736
rect 5648 8676 5652 8732
rect 5652 8676 5708 8732
rect 5708 8676 5712 8732
rect 5648 8672 5712 8676
rect 5728 8732 5792 8736
rect 5728 8676 5732 8732
rect 5732 8676 5788 8732
rect 5788 8676 5792 8732
rect 5728 8672 5792 8676
rect 5808 8732 5872 8736
rect 5808 8676 5812 8732
rect 5812 8676 5868 8732
rect 5868 8676 5872 8732
rect 5808 8672 5872 8676
rect 5888 8732 5952 8736
rect 5888 8676 5892 8732
rect 5892 8676 5948 8732
rect 5948 8676 5952 8732
rect 5888 8672 5952 8676
rect 8339 8732 8403 8736
rect 8339 8676 8343 8732
rect 8343 8676 8399 8732
rect 8399 8676 8403 8732
rect 8339 8672 8403 8676
rect 8419 8732 8483 8736
rect 8419 8676 8423 8732
rect 8423 8676 8479 8732
rect 8479 8676 8483 8732
rect 8419 8672 8483 8676
rect 8499 8732 8563 8736
rect 8499 8676 8503 8732
rect 8503 8676 8559 8732
rect 8559 8676 8563 8732
rect 8499 8672 8563 8676
rect 8579 8732 8643 8736
rect 8579 8676 8583 8732
rect 8583 8676 8639 8732
rect 8639 8676 8643 8732
rect 8579 8672 8643 8676
rect 11030 8732 11094 8736
rect 11030 8676 11034 8732
rect 11034 8676 11090 8732
rect 11090 8676 11094 8732
rect 11030 8672 11094 8676
rect 11110 8732 11174 8736
rect 11110 8676 11114 8732
rect 11114 8676 11170 8732
rect 11170 8676 11174 8732
rect 11110 8672 11174 8676
rect 11190 8732 11254 8736
rect 11190 8676 11194 8732
rect 11194 8676 11250 8732
rect 11250 8676 11254 8732
rect 11190 8672 11254 8676
rect 11270 8732 11334 8736
rect 11270 8676 11274 8732
rect 11274 8676 11330 8732
rect 11330 8676 11334 8732
rect 11270 8672 11334 8676
rect 2297 8188 2361 8192
rect 2297 8132 2301 8188
rect 2301 8132 2357 8188
rect 2357 8132 2361 8188
rect 2297 8128 2361 8132
rect 2377 8188 2441 8192
rect 2377 8132 2381 8188
rect 2381 8132 2437 8188
rect 2437 8132 2441 8188
rect 2377 8128 2441 8132
rect 2457 8188 2521 8192
rect 2457 8132 2461 8188
rect 2461 8132 2517 8188
rect 2517 8132 2521 8188
rect 2457 8128 2521 8132
rect 2537 8188 2601 8192
rect 2537 8132 2541 8188
rect 2541 8132 2597 8188
rect 2597 8132 2601 8188
rect 2537 8128 2601 8132
rect 4988 8188 5052 8192
rect 4988 8132 4992 8188
rect 4992 8132 5048 8188
rect 5048 8132 5052 8188
rect 4988 8128 5052 8132
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 7679 8188 7743 8192
rect 7679 8132 7683 8188
rect 7683 8132 7739 8188
rect 7739 8132 7743 8188
rect 7679 8128 7743 8132
rect 7759 8188 7823 8192
rect 7759 8132 7763 8188
rect 7763 8132 7819 8188
rect 7819 8132 7823 8188
rect 7759 8128 7823 8132
rect 7839 8188 7903 8192
rect 7839 8132 7843 8188
rect 7843 8132 7899 8188
rect 7899 8132 7903 8188
rect 7839 8128 7903 8132
rect 7919 8188 7983 8192
rect 7919 8132 7923 8188
rect 7923 8132 7979 8188
rect 7979 8132 7983 8188
rect 7919 8128 7983 8132
rect 10370 8188 10434 8192
rect 10370 8132 10374 8188
rect 10374 8132 10430 8188
rect 10430 8132 10434 8188
rect 10370 8128 10434 8132
rect 10450 8188 10514 8192
rect 10450 8132 10454 8188
rect 10454 8132 10510 8188
rect 10510 8132 10514 8188
rect 10450 8128 10514 8132
rect 10530 8188 10594 8192
rect 10530 8132 10534 8188
rect 10534 8132 10590 8188
rect 10590 8132 10594 8188
rect 10530 8128 10594 8132
rect 10610 8188 10674 8192
rect 10610 8132 10614 8188
rect 10614 8132 10670 8188
rect 10670 8132 10674 8188
rect 10610 8128 10674 8132
rect 2957 7644 3021 7648
rect 2957 7588 2961 7644
rect 2961 7588 3017 7644
rect 3017 7588 3021 7644
rect 2957 7584 3021 7588
rect 3037 7644 3101 7648
rect 3037 7588 3041 7644
rect 3041 7588 3097 7644
rect 3097 7588 3101 7644
rect 3037 7584 3101 7588
rect 3117 7644 3181 7648
rect 3117 7588 3121 7644
rect 3121 7588 3177 7644
rect 3177 7588 3181 7644
rect 3117 7584 3181 7588
rect 3197 7644 3261 7648
rect 3197 7588 3201 7644
rect 3201 7588 3257 7644
rect 3257 7588 3261 7644
rect 3197 7584 3261 7588
rect 5648 7644 5712 7648
rect 5648 7588 5652 7644
rect 5652 7588 5708 7644
rect 5708 7588 5712 7644
rect 5648 7584 5712 7588
rect 5728 7644 5792 7648
rect 5728 7588 5732 7644
rect 5732 7588 5788 7644
rect 5788 7588 5792 7644
rect 5728 7584 5792 7588
rect 5808 7644 5872 7648
rect 5808 7588 5812 7644
rect 5812 7588 5868 7644
rect 5868 7588 5872 7644
rect 5808 7584 5872 7588
rect 5888 7644 5952 7648
rect 5888 7588 5892 7644
rect 5892 7588 5948 7644
rect 5948 7588 5952 7644
rect 5888 7584 5952 7588
rect 8339 7644 8403 7648
rect 8339 7588 8343 7644
rect 8343 7588 8399 7644
rect 8399 7588 8403 7644
rect 8339 7584 8403 7588
rect 8419 7644 8483 7648
rect 8419 7588 8423 7644
rect 8423 7588 8479 7644
rect 8479 7588 8483 7644
rect 8419 7584 8483 7588
rect 8499 7644 8563 7648
rect 8499 7588 8503 7644
rect 8503 7588 8559 7644
rect 8559 7588 8563 7644
rect 8499 7584 8563 7588
rect 8579 7644 8643 7648
rect 8579 7588 8583 7644
rect 8583 7588 8639 7644
rect 8639 7588 8643 7644
rect 8579 7584 8643 7588
rect 11030 7644 11094 7648
rect 11030 7588 11034 7644
rect 11034 7588 11090 7644
rect 11090 7588 11094 7644
rect 11030 7584 11094 7588
rect 11110 7644 11174 7648
rect 11110 7588 11114 7644
rect 11114 7588 11170 7644
rect 11170 7588 11174 7644
rect 11110 7584 11174 7588
rect 11190 7644 11254 7648
rect 11190 7588 11194 7644
rect 11194 7588 11250 7644
rect 11250 7588 11254 7644
rect 11190 7584 11254 7588
rect 11270 7644 11334 7648
rect 11270 7588 11274 7644
rect 11274 7588 11330 7644
rect 11330 7588 11334 7644
rect 11270 7584 11334 7588
rect 2297 7100 2361 7104
rect 2297 7044 2301 7100
rect 2301 7044 2357 7100
rect 2357 7044 2361 7100
rect 2297 7040 2361 7044
rect 2377 7100 2441 7104
rect 2377 7044 2381 7100
rect 2381 7044 2437 7100
rect 2437 7044 2441 7100
rect 2377 7040 2441 7044
rect 2457 7100 2521 7104
rect 2457 7044 2461 7100
rect 2461 7044 2517 7100
rect 2517 7044 2521 7100
rect 2457 7040 2521 7044
rect 2537 7100 2601 7104
rect 2537 7044 2541 7100
rect 2541 7044 2597 7100
rect 2597 7044 2601 7100
rect 2537 7040 2601 7044
rect 4988 7100 5052 7104
rect 4988 7044 4992 7100
rect 4992 7044 5048 7100
rect 5048 7044 5052 7100
rect 4988 7040 5052 7044
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 7679 7100 7743 7104
rect 7679 7044 7683 7100
rect 7683 7044 7739 7100
rect 7739 7044 7743 7100
rect 7679 7040 7743 7044
rect 7759 7100 7823 7104
rect 7759 7044 7763 7100
rect 7763 7044 7819 7100
rect 7819 7044 7823 7100
rect 7759 7040 7823 7044
rect 7839 7100 7903 7104
rect 7839 7044 7843 7100
rect 7843 7044 7899 7100
rect 7899 7044 7903 7100
rect 7839 7040 7903 7044
rect 7919 7100 7983 7104
rect 7919 7044 7923 7100
rect 7923 7044 7979 7100
rect 7979 7044 7983 7100
rect 7919 7040 7983 7044
rect 10370 7100 10434 7104
rect 10370 7044 10374 7100
rect 10374 7044 10430 7100
rect 10430 7044 10434 7100
rect 10370 7040 10434 7044
rect 10450 7100 10514 7104
rect 10450 7044 10454 7100
rect 10454 7044 10510 7100
rect 10510 7044 10514 7100
rect 10450 7040 10514 7044
rect 10530 7100 10594 7104
rect 10530 7044 10534 7100
rect 10534 7044 10590 7100
rect 10590 7044 10594 7100
rect 10530 7040 10594 7044
rect 10610 7100 10674 7104
rect 10610 7044 10614 7100
rect 10614 7044 10670 7100
rect 10670 7044 10674 7100
rect 10610 7040 10674 7044
rect 2957 6556 3021 6560
rect 2957 6500 2961 6556
rect 2961 6500 3017 6556
rect 3017 6500 3021 6556
rect 2957 6496 3021 6500
rect 3037 6556 3101 6560
rect 3037 6500 3041 6556
rect 3041 6500 3097 6556
rect 3097 6500 3101 6556
rect 3037 6496 3101 6500
rect 3117 6556 3181 6560
rect 3117 6500 3121 6556
rect 3121 6500 3177 6556
rect 3177 6500 3181 6556
rect 3117 6496 3181 6500
rect 3197 6556 3261 6560
rect 3197 6500 3201 6556
rect 3201 6500 3257 6556
rect 3257 6500 3261 6556
rect 3197 6496 3261 6500
rect 5648 6556 5712 6560
rect 5648 6500 5652 6556
rect 5652 6500 5708 6556
rect 5708 6500 5712 6556
rect 5648 6496 5712 6500
rect 5728 6556 5792 6560
rect 5728 6500 5732 6556
rect 5732 6500 5788 6556
rect 5788 6500 5792 6556
rect 5728 6496 5792 6500
rect 5808 6556 5872 6560
rect 5808 6500 5812 6556
rect 5812 6500 5868 6556
rect 5868 6500 5872 6556
rect 5808 6496 5872 6500
rect 5888 6556 5952 6560
rect 5888 6500 5892 6556
rect 5892 6500 5948 6556
rect 5948 6500 5952 6556
rect 5888 6496 5952 6500
rect 8339 6556 8403 6560
rect 8339 6500 8343 6556
rect 8343 6500 8399 6556
rect 8399 6500 8403 6556
rect 8339 6496 8403 6500
rect 8419 6556 8483 6560
rect 8419 6500 8423 6556
rect 8423 6500 8479 6556
rect 8479 6500 8483 6556
rect 8419 6496 8483 6500
rect 8499 6556 8563 6560
rect 8499 6500 8503 6556
rect 8503 6500 8559 6556
rect 8559 6500 8563 6556
rect 8499 6496 8563 6500
rect 8579 6556 8643 6560
rect 8579 6500 8583 6556
rect 8583 6500 8639 6556
rect 8639 6500 8643 6556
rect 8579 6496 8643 6500
rect 11030 6556 11094 6560
rect 11030 6500 11034 6556
rect 11034 6500 11090 6556
rect 11090 6500 11094 6556
rect 11030 6496 11094 6500
rect 11110 6556 11174 6560
rect 11110 6500 11114 6556
rect 11114 6500 11170 6556
rect 11170 6500 11174 6556
rect 11110 6496 11174 6500
rect 11190 6556 11254 6560
rect 11190 6500 11194 6556
rect 11194 6500 11250 6556
rect 11250 6500 11254 6556
rect 11190 6496 11254 6500
rect 11270 6556 11334 6560
rect 11270 6500 11274 6556
rect 11274 6500 11330 6556
rect 11330 6500 11334 6556
rect 11270 6496 11334 6500
rect 2297 6012 2361 6016
rect 2297 5956 2301 6012
rect 2301 5956 2357 6012
rect 2357 5956 2361 6012
rect 2297 5952 2361 5956
rect 2377 6012 2441 6016
rect 2377 5956 2381 6012
rect 2381 5956 2437 6012
rect 2437 5956 2441 6012
rect 2377 5952 2441 5956
rect 2457 6012 2521 6016
rect 2457 5956 2461 6012
rect 2461 5956 2517 6012
rect 2517 5956 2521 6012
rect 2457 5952 2521 5956
rect 2537 6012 2601 6016
rect 2537 5956 2541 6012
rect 2541 5956 2597 6012
rect 2597 5956 2601 6012
rect 2537 5952 2601 5956
rect 4988 6012 5052 6016
rect 4988 5956 4992 6012
rect 4992 5956 5048 6012
rect 5048 5956 5052 6012
rect 4988 5952 5052 5956
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 7679 6012 7743 6016
rect 7679 5956 7683 6012
rect 7683 5956 7739 6012
rect 7739 5956 7743 6012
rect 7679 5952 7743 5956
rect 7759 6012 7823 6016
rect 7759 5956 7763 6012
rect 7763 5956 7819 6012
rect 7819 5956 7823 6012
rect 7759 5952 7823 5956
rect 7839 6012 7903 6016
rect 7839 5956 7843 6012
rect 7843 5956 7899 6012
rect 7899 5956 7903 6012
rect 7839 5952 7903 5956
rect 7919 6012 7983 6016
rect 7919 5956 7923 6012
rect 7923 5956 7979 6012
rect 7979 5956 7983 6012
rect 7919 5952 7983 5956
rect 10370 6012 10434 6016
rect 10370 5956 10374 6012
rect 10374 5956 10430 6012
rect 10430 5956 10434 6012
rect 10370 5952 10434 5956
rect 10450 6012 10514 6016
rect 10450 5956 10454 6012
rect 10454 5956 10510 6012
rect 10510 5956 10514 6012
rect 10450 5952 10514 5956
rect 10530 6012 10594 6016
rect 10530 5956 10534 6012
rect 10534 5956 10590 6012
rect 10590 5956 10594 6012
rect 10530 5952 10594 5956
rect 10610 6012 10674 6016
rect 10610 5956 10614 6012
rect 10614 5956 10670 6012
rect 10670 5956 10674 6012
rect 10610 5952 10674 5956
rect 2957 5468 3021 5472
rect 2957 5412 2961 5468
rect 2961 5412 3017 5468
rect 3017 5412 3021 5468
rect 2957 5408 3021 5412
rect 3037 5468 3101 5472
rect 3037 5412 3041 5468
rect 3041 5412 3097 5468
rect 3097 5412 3101 5468
rect 3037 5408 3101 5412
rect 3117 5468 3181 5472
rect 3117 5412 3121 5468
rect 3121 5412 3177 5468
rect 3177 5412 3181 5468
rect 3117 5408 3181 5412
rect 3197 5468 3261 5472
rect 3197 5412 3201 5468
rect 3201 5412 3257 5468
rect 3257 5412 3261 5468
rect 3197 5408 3261 5412
rect 5648 5468 5712 5472
rect 5648 5412 5652 5468
rect 5652 5412 5708 5468
rect 5708 5412 5712 5468
rect 5648 5408 5712 5412
rect 5728 5468 5792 5472
rect 5728 5412 5732 5468
rect 5732 5412 5788 5468
rect 5788 5412 5792 5468
rect 5728 5408 5792 5412
rect 5808 5468 5872 5472
rect 5808 5412 5812 5468
rect 5812 5412 5868 5468
rect 5868 5412 5872 5468
rect 5808 5408 5872 5412
rect 5888 5468 5952 5472
rect 5888 5412 5892 5468
rect 5892 5412 5948 5468
rect 5948 5412 5952 5468
rect 5888 5408 5952 5412
rect 8339 5468 8403 5472
rect 8339 5412 8343 5468
rect 8343 5412 8399 5468
rect 8399 5412 8403 5468
rect 8339 5408 8403 5412
rect 8419 5468 8483 5472
rect 8419 5412 8423 5468
rect 8423 5412 8479 5468
rect 8479 5412 8483 5468
rect 8419 5408 8483 5412
rect 8499 5468 8563 5472
rect 8499 5412 8503 5468
rect 8503 5412 8559 5468
rect 8559 5412 8563 5468
rect 8499 5408 8563 5412
rect 8579 5468 8643 5472
rect 8579 5412 8583 5468
rect 8583 5412 8639 5468
rect 8639 5412 8643 5468
rect 8579 5408 8643 5412
rect 11030 5468 11094 5472
rect 11030 5412 11034 5468
rect 11034 5412 11090 5468
rect 11090 5412 11094 5468
rect 11030 5408 11094 5412
rect 11110 5468 11174 5472
rect 11110 5412 11114 5468
rect 11114 5412 11170 5468
rect 11170 5412 11174 5468
rect 11110 5408 11174 5412
rect 11190 5468 11254 5472
rect 11190 5412 11194 5468
rect 11194 5412 11250 5468
rect 11250 5412 11254 5468
rect 11190 5408 11254 5412
rect 11270 5468 11334 5472
rect 11270 5412 11274 5468
rect 11274 5412 11330 5468
rect 11330 5412 11334 5468
rect 11270 5408 11334 5412
rect 2297 4924 2361 4928
rect 2297 4868 2301 4924
rect 2301 4868 2357 4924
rect 2357 4868 2361 4924
rect 2297 4864 2361 4868
rect 2377 4924 2441 4928
rect 2377 4868 2381 4924
rect 2381 4868 2437 4924
rect 2437 4868 2441 4924
rect 2377 4864 2441 4868
rect 2457 4924 2521 4928
rect 2457 4868 2461 4924
rect 2461 4868 2517 4924
rect 2517 4868 2521 4924
rect 2457 4864 2521 4868
rect 2537 4924 2601 4928
rect 2537 4868 2541 4924
rect 2541 4868 2597 4924
rect 2597 4868 2601 4924
rect 2537 4864 2601 4868
rect 4988 4924 5052 4928
rect 4988 4868 4992 4924
rect 4992 4868 5048 4924
rect 5048 4868 5052 4924
rect 4988 4864 5052 4868
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 7679 4924 7743 4928
rect 7679 4868 7683 4924
rect 7683 4868 7739 4924
rect 7739 4868 7743 4924
rect 7679 4864 7743 4868
rect 7759 4924 7823 4928
rect 7759 4868 7763 4924
rect 7763 4868 7819 4924
rect 7819 4868 7823 4924
rect 7759 4864 7823 4868
rect 7839 4924 7903 4928
rect 7839 4868 7843 4924
rect 7843 4868 7899 4924
rect 7899 4868 7903 4924
rect 7839 4864 7903 4868
rect 7919 4924 7983 4928
rect 7919 4868 7923 4924
rect 7923 4868 7979 4924
rect 7979 4868 7983 4924
rect 7919 4864 7983 4868
rect 10370 4924 10434 4928
rect 10370 4868 10374 4924
rect 10374 4868 10430 4924
rect 10430 4868 10434 4924
rect 10370 4864 10434 4868
rect 10450 4924 10514 4928
rect 10450 4868 10454 4924
rect 10454 4868 10510 4924
rect 10510 4868 10514 4924
rect 10450 4864 10514 4868
rect 10530 4924 10594 4928
rect 10530 4868 10534 4924
rect 10534 4868 10590 4924
rect 10590 4868 10594 4924
rect 10530 4864 10594 4868
rect 10610 4924 10674 4928
rect 10610 4868 10614 4924
rect 10614 4868 10670 4924
rect 10670 4868 10674 4924
rect 10610 4864 10674 4868
rect 2957 4380 3021 4384
rect 2957 4324 2961 4380
rect 2961 4324 3017 4380
rect 3017 4324 3021 4380
rect 2957 4320 3021 4324
rect 3037 4380 3101 4384
rect 3037 4324 3041 4380
rect 3041 4324 3097 4380
rect 3097 4324 3101 4380
rect 3037 4320 3101 4324
rect 3117 4380 3181 4384
rect 3117 4324 3121 4380
rect 3121 4324 3177 4380
rect 3177 4324 3181 4380
rect 3117 4320 3181 4324
rect 3197 4380 3261 4384
rect 3197 4324 3201 4380
rect 3201 4324 3257 4380
rect 3257 4324 3261 4380
rect 3197 4320 3261 4324
rect 5648 4380 5712 4384
rect 5648 4324 5652 4380
rect 5652 4324 5708 4380
rect 5708 4324 5712 4380
rect 5648 4320 5712 4324
rect 5728 4380 5792 4384
rect 5728 4324 5732 4380
rect 5732 4324 5788 4380
rect 5788 4324 5792 4380
rect 5728 4320 5792 4324
rect 5808 4380 5872 4384
rect 5808 4324 5812 4380
rect 5812 4324 5868 4380
rect 5868 4324 5872 4380
rect 5808 4320 5872 4324
rect 5888 4380 5952 4384
rect 5888 4324 5892 4380
rect 5892 4324 5948 4380
rect 5948 4324 5952 4380
rect 5888 4320 5952 4324
rect 8339 4380 8403 4384
rect 8339 4324 8343 4380
rect 8343 4324 8399 4380
rect 8399 4324 8403 4380
rect 8339 4320 8403 4324
rect 8419 4380 8483 4384
rect 8419 4324 8423 4380
rect 8423 4324 8479 4380
rect 8479 4324 8483 4380
rect 8419 4320 8483 4324
rect 8499 4380 8563 4384
rect 8499 4324 8503 4380
rect 8503 4324 8559 4380
rect 8559 4324 8563 4380
rect 8499 4320 8563 4324
rect 8579 4380 8643 4384
rect 8579 4324 8583 4380
rect 8583 4324 8639 4380
rect 8639 4324 8643 4380
rect 8579 4320 8643 4324
rect 11030 4380 11094 4384
rect 11030 4324 11034 4380
rect 11034 4324 11090 4380
rect 11090 4324 11094 4380
rect 11030 4320 11094 4324
rect 11110 4380 11174 4384
rect 11110 4324 11114 4380
rect 11114 4324 11170 4380
rect 11170 4324 11174 4380
rect 11110 4320 11174 4324
rect 11190 4380 11254 4384
rect 11190 4324 11194 4380
rect 11194 4324 11250 4380
rect 11250 4324 11254 4380
rect 11190 4320 11254 4324
rect 11270 4380 11334 4384
rect 11270 4324 11274 4380
rect 11274 4324 11330 4380
rect 11330 4324 11334 4380
rect 11270 4320 11334 4324
rect 2297 3836 2361 3840
rect 2297 3780 2301 3836
rect 2301 3780 2357 3836
rect 2357 3780 2361 3836
rect 2297 3776 2361 3780
rect 2377 3836 2441 3840
rect 2377 3780 2381 3836
rect 2381 3780 2437 3836
rect 2437 3780 2441 3836
rect 2377 3776 2441 3780
rect 2457 3836 2521 3840
rect 2457 3780 2461 3836
rect 2461 3780 2517 3836
rect 2517 3780 2521 3836
rect 2457 3776 2521 3780
rect 2537 3836 2601 3840
rect 2537 3780 2541 3836
rect 2541 3780 2597 3836
rect 2597 3780 2601 3836
rect 2537 3776 2601 3780
rect 4988 3836 5052 3840
rect 4988 3780 4992 3836
rect 4992 3780 5048 3836
rect 5048 3780 5052 3836
rect 4988 3776 5052 3780
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 7679 3836 7743 3840
rect 7679 3780 7683 3836
rect 7683 3780 7739 3836
rect 7739 3780 7743 3836
rect 7679 3776 7743 3780
rect 7759 3836 7823 3840
rect 7759 3780 7763 3836
rect 7763 3780 7819 3836
rect 7819 3780 7823 3836
rect 7759 3776 7823 3780
rect 7839 3836 7903 3840
rect 7839 3780 7843 3836
rect 7843 3780 7899 3836
rect 7899 3780 7903 3836
rect 7839 3776 7903 3780
rect 7919 3836 7983 3840
rect 7919 3780 7923 3836
rect 7923 3780 7979 3836
rect 7979 3780 7983 3836
rect 7919 3776 7983 3780
rect 10370 3836 10434 3840
rect 10370 3780 10374 3836
rect 10374 3780 10430 3836
rect 10430 3780 10434 3836
rect 10370 3776 10434 3780
rect 10450 3836 10514 3840
rect 10450 3780 10454 3836
rect 10454 3780 10510 3836
rect 10510 3780 10514 3836
rect 10450 3776 10514 3780
rect 10530 3836 10594 3840
rect 10530 3780 10534 3836
rect 10534 3780 10590 3836
rect 10590 3780 10594 3836
rect 10530 3776 10594 3780
rect 10610 3836 10674 3840
rect 10610 3780 10614 3836
rect 10614 3780 10670 3836
rect 10670 3780 10674 3836
rect 10610 3776 10674 3780
rect 2957 3292 3021 3296
rect 2957 3236 2961 3292
rect 2961 3236 3017 3292
rect 3017 3236 3021 3292
rect 2957 3232 3021 3236
rect 3037 3292 3101 3296
rect 3037 3236 3041 3292
rect 3041 3236 3097 3292
rect 3097 3236 3101 3292
rect 3037 3232 3101 3236
rect 3117 3292 3181 3296
rect 3117 3236 3121 3292
rect 3121 3236 3177 3292
rect 3177 3236 3181 3292
rect 3117 3232 3181 3236
rect 3197 3292 3261 3296
rect 3197 3236 3201 3292
rect 3201 3236 3257 3292
rect 3257 3236 3261 3292
rect 3197 3232 3261 3236
rect 5648 3292 5712 3296
rect 5648 3236 5652 3292
rect 5652 3236 5708 3292
rect 5708 3236 5712 3292
rect 5648 3232 5712 3236
rect 5728 3292 5792 3296
rect 5728 3236 5732 3292
rect 5732 3236 5788 3292
rect 5788 3236 5792 3292
rect 5728 3232 5792 3236
rect 5808 3292 5872 3296
rect 5808 3236 5812 3292
rect 5812 3236 5868 3292
rect 5868 3236 5872 3292
rect 5808 3232 5872 3236
rect 5888 3292 5952 3296
rect 5888 3236 5892 3292
rect 5892 3236 5948 3292
rect 5948 3236 5952 3292
rect 5888 3232 5952 3236
rect 8339 3292 8403 3296
rect 8339 3236 8343 3292
rect 8343 3236 8399 3292
rect 8399 3236 8403 3292
rect 8339 3232 8403 3236
rect 8419 3292 8483 3296
rect 8419 3236 8423 3292
rect 8423 3236 8479 3292
rect 8479 3236 8483 3292
rect 8419 3232 8483 3236
rect 8499 3292 8563 3296
rect 8499 3236 8503 3292
rect 8503 3236 8559 3292
rect 8559 3236 8563 3292
rect 8499 3232 8563 3236
rect 8579 3292 8643 3296
rect 8579 3236 8583 3292
rect 8583 3236 8639 3292
rect 8639 3236 8643 3292
rect 8579 3232 8643 3236
rect 11030 3292 11094 3296
rect 11030 3236 11034 3292
rect 11034 3236 11090 3292
rect 11090 3236 11094 3292
rect 11030 3232 11094 3236
rect 11110 3292 11174 3296
rect 11110 3236 11114 3292
rect 11114 3236 11170 3292
rect 11170 3236 11174 3292
rect 11110 3232 11174 3236
rect 11190 3292 11254 3296
rect 11190 3236 11194 3292
rect 11194 3236 11250 3292
rect 11250 3236 11254 3292
rect 11190 3232 11254 3236
rect 11270 3292 11334 3296
rect 11270 3236 11274 3292
rect 11274 3236 11330 3292
rect 11330 3236 11334 3292
rect 11270 3232 11334 3236
rect 2297 2748 2361 2752
rect 2297 2692 2301 2748
rect 2301 2692 2357 2748
rect 2357 2692 2361 2748
rect 2297 2688 2361 2692
rect 2377 2748 2441 2752
rect 2377 2692 2381 2748
rect 2381 2692 2437 2748
rect 2437 2692 2441 2748
rect 2377 2688 2441 2692
rect 2457 2748 2521 2752
rect 2457 2692 2461 2748
rect 2461 2692 2517 2748
rect 2517 2692 2521 2748
rect 2457 2688 2521 2692
rect 2537 2748 2601 2752
rect 2537 2692 2541 2748
rect 2541 2692 2597 2748
rect 2597 2692 2601 2748
rect 2537 2688 2601 2692
rect 4988 2748 5052 2752
rect 4988 2692 4992 2748
rect 4992 2692 5048 2748
rect 5048 2692 5052 2748
rect 4988 2688 5052 2692
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 7679 2748 7743 2752
rect 7679 2692 7683 2748
rect 7683 2692 7739 2748
rect 7739 2692 7743 2748
rect 7679 2688 7743 2692
rect 7759 2748 7823 2752
rect 7759 2692 7763 2748
rect 7763 2692 7819 2748
rect 7819 2692 7823 2748
rect 7759 2688 7823 2692
rect 7839 2748 7903 2752
rect 7839 2692 7843 2748
rect 7843 2692 7899 2748
rect 7899 2692 7903 2748
rect 7839 2688 7903 2692
rect 7919 2748 7983 2752
rect 7919 2692 7923 2748
rect 7923 2692 7979 2748
rect 7979 2692 7983 2748
rect 7919 2688 7983 2692
rect 10370 2748 10434 2752
rect 10370 2692 10374 2748
rect 10374 2692 10430 2748
rect 10430 2692 10434 2748
rect 10370 2688 10434 2692
rect 10450 2748 10514 2752
rect 10450 2692 10454 2748
rect 10454 2692 10510 2748
rect 10510 2692 10514 2748
rect 10450 2688 10514 2692
rect 10530 2748 10594 2752
rect 10530 2692 10534 2748
rect 10534 2692 10590 2748
rect 10590 2692 10594 2748
rect 10530 2688 10594 2692
rect 10610 2748 10674 2752
rect 10610 2692 10614 2748
rect 10614 2692 10670 2748
rect 10670 2692 10674 2748
rect 10610 2688 10674 2692
rect 7420 2680 7484 2684
rect 7420 2624 7470 2680
rect 7470 2624 7484 2680
rect 7420 2620 7484 2624
rect 2957 2204 3021 2208
rect 2957 2148 2961 2204
rect 2961 2148 3017 2204
rect 3017 2148 3021 2204
rect 2957 2144 3021 2148
rect 3037 2204 3101 2208
rect 3037 2148 3041 2204
rect 3041 2148 3097 2204
rect 3097 2148 3101 2204
rect 3037 2144 3101 2148
rect 3117 2204 3181 2208
rect 3117 2148 3121 2204
rect 3121 2148 3177 2204
rect 3177 2148 3181 2204
rect 3117 2144 3181 2148
rect 3197 2204 3261 2208
rect 3197 2148 3201 2204
rect 3201 2148 3257 2204
rect 3257 2148 3261 2204
rect 3197 2144 3261 2148
rect 5648 2204 5712 2208
rect 5648 2148 5652 2204
rect 5652 2148 5708 2204
rect 5708 2148 5712 2204
rect 5648 2144 5712 2148
rect 5728 2204 5792 2208
rect 5728 2148 5732 2204
rect 5732 2148 5788 2204
rect 5788 2148 5792 2204
rect 5728 2144 5792 2148
rect 5808 2204 5872 2208
rect 5808 2148 5812 2204
rect 5812 2148 5868 2204
rect 5868 2148 5872 2204
rect 5808 2144 5872 2148
rect 5888 2204 5952 2208
rect 5888 2148 5892 2204
rect 5892 2148 5948 2204
rect 5948 2148 5952 2204
rect 5888 2144 5952 2148
rect 8339 2204 8403 2208
rect 8339 2148 8343 2204
rect 8343 2148 8399 2204
rect 8399 2148 8403 2204
rect 8339 2144 8403 2148
rect 8419 2204 8483 2208
rect 8419 2148 8423 2204
rect 8423 2148 8479 2204
rect 8479 2148 8483 2204
rect 8419 2144 8483 2148
rect 8499 2204 8563 2208
rect 8499 2148 8503 2204
rect 8503 2148 8559 2204
rect 8559 2148 8563 2204
rect 8499 2144 8563 2148
rect 8579 2204 8643 2208
rect 8579 2148 8583 2204
rect 8583 2148 8639 2204
rect 8639 2148 8643 2204
rect 8579 2144 8643 2148
rect 11030 2204 11094 2208
rect 11030 2148 11034 2204
rect 11034 2148 11090 2204
rect 11090 2148 11094 2204
rect 11030 2144 11094 2148
rect 11110 2204 11174 2208
rect 11110 2148 11114 2204
rect 11114 2148 11170 2204
rect 11170 2148 11174 2204
rect 11110 2144 11174 2148
rect 11190 2204 11254 2208
rect 11190 2148 11194 2204
rect 11194 2148 11250 2204
rect 11250 2148 11254 2204
rect 11190 2144 11254 2148
rect 11270 2204 11334 2208
rect 11270 2148 11274 2204
rect 11274 2148 11330 2204
rect 11330 2148 11334 2204
rect 11270 2144 11334 2148
<< metal4 >>
rect 2289 12544 2609 12560
rect 2289 12480 2297 12544
rect 2361 12480 2377 12544
rect 2441 12480 2457 12544
rect 2521 12480 2537 12544
rect 2601 12480 2609 12544
rect 2289 11456 2609 12480
rect 2289 11392 2297 11456
rect 2361 11392 2377 11456
rect 2441 11392 2457 11456
rect 2521 11392 2537 11456
rect 2601 11392 2609 11456
rect 2289 11338 2609 11392
rect 2289 11102 2331 11338
rect 2567 11102 2609 11338
rect 2289 10368 2609 11102
rect 2289 10304 2297 10368
rect 2361 10304 2377 10368
rect 2441 10304 2457 10368
rect 2521 10304 2537 10368
rect 2601 10304 2609 10368
rect 2289 9280 2609 10304
rect 2289 9216 2297 9280
rect 2361 9216 2377 9280
rect 2441 9216 2457 9280
rect 2521 9216 2537 9280
rect 2601 9216 2609 9280
rect 2289 8754 2609 9216
rect 2289 8518 2331 8754
rect 2567 8518 2609 8754
rect 2289 8192 2609 8518
rect 2289 8128 2297 8192
rect 2361 8128 2377 8192
rect 2441 8128 2457 8192
rect 2521 8128 2537 8192
rect 2601 8128 2609 8192
rect 2289 7104 2609 8128
rect 2289 7040 2297 7104
rect 2361 7040 2377 7104
rect 2441 7040 2457 7104
rect 2521 7040 2537 7104
rect 2601 7040 2609 7104
rect 2289 6170 2609 7040
rect 2289 6016 2331 6170
rect 2567 6016 2609 6170
rect 2289 5952 2297 6016
rect 2601 5952 2609 6016
rect 2289 5934 2331 5952
rect 2567 5934 2609 5952
rect 2289 4928 2609 5934
rect 2289 4864 2297 4928
rect 2361 4864 2377 4928
rect 2441 4864 2457 4928
rect 2521 4864 2537 4928
rect 2601 4864 2609 4928
rect 2289 3840 2609 4864
rect 2289 3776 2297 3840
rect 2361 3776 2377 3840
rect 2441 3776 2457 3840
rect 2521 3776 2537 3840
rect 2601 3776 2609 3840
rect 2289 3586 2609 3776
rect 2289 3350 2331 3586
rect 2567 3350 2609 3586
rect 2289 2752 2609 3350
rect 2289 2688 2297 2752
rect 2361 2688 2377 2752
rect 2441 2688 2457 2752
rect 2521 2688 2537 2752
rect 2601 2688 2609 2752
rect 2289 2128 2609 2688
rect 2949 12000 3269 12560
rect 2949 11936 2957 12000
rect 3021 11998 3037 12000
rect 3101 11998 3117 12000
rect 3181 11998 3197 12000
rect 3261 11936 3269 12000
rect 2949 11762 2991 11936
rect 3227 11762 3269 11936
rect 2949 10912 3269 11762
rect 2949 10848 2957 10912
rect 3021 10848 3037 10912
rect 3101 10848 3117 10912
rect 3181 10848 3197 10912
rect 3261 10848 3269 10912
rect 2949 9824 3269 10848
rect 2949 9760 2957 9824
rect 3021 9760 3037 9824
rect 3101 9760 3117 9824
rect 3181 9760 3197 9824
rect 3261 9760 3269 9824
rect 2949 9414 3269 9760
rect 2949 9178 2991 9414
rect 3227 9178 3269 9414
rect 2949 8736 3269 9178
rect 2949 8672 2957 8736
rect 3021 8672 3037 8736
rect 3101 8672 3117 8736
rect 3181 8672 3197 8736
rect 3261 8672 3269 8736
rect 2949 7648 3269 8672
rect 2949 7584 2957 7648
rect 3021 7584 3037 7648
rect 3101 7584 3117 7648
rect 3181 7584 3197 7648
rect 3261 7584 3269 7648
rect 2949 6830 3269 7584
rect 2949 6594 2991 6830
rect 3227 6594 3269 6830
rect 2949 6560 3269 6594
rect 2949 6496 2957 6560
rect 3021 6496 3037 6560
rect 3101 6496 3117 6560
rect 3181 6496 3197 6560
rect 3261 6496 3269 6560
rect 2949 5472 3269 6496
rect 2949 5408 2957 5472
rect 3021 5408 3037 5472
rect 3101 5408 3117 5472
rect 3181 5408 3197 5472
rect 3261 5408 3269 5472
rect 2949 4384 3269 5408
rect 2949 4320 2957 4384
rect 3021 4320 3037 4384
rect 3101 4320 3117 4384
rect 3181 4320 3197 4384
rect 3261 4320 3269 4384
rect 2949 4246 3269 4320
rect 2949 4010 2991 4246
rect 3227 4010 3269 4246
rect 2949 3296 3269 4010
rect 2949 3232 2957 3296
rect 3021 3232 3037 3296
rect 3101 3232 3117 3296
rect 3181 3232 3197 3296
rect 3261 3232 3269 3296
rect 2949 2208 3269 3232
rect 2949 2144 2957 2208
rect 3021 2144 3037 2208
rect 3101 2144 3117 2208
rect 3181 2144 3197 2208
rect 3261 2144 3269 2208
rect 2949 2128 3269 2144
rect 4980 12544 5300 12560
rect 4980 12480 4988 12544
rect 5052 12480 5068 12544
rect 5132 12480 5148 12544
rect 5212 12480 5228 12544
rect 5292 12480 5300 12544
rect 4980 11456 5300 12480
rect 4980 11392 4988 11456
rect 5052 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5300 11456
rect 4980 11338 5300 11392
rect 4980 11102 5022 11338
rect 5258 11102 5300 11338
rect 4980 10368 5300 11102
rect 4980 10304 4988 10368
rect 5052 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5300 10368
rect 4980 9280 5300 10304
rect 4980 9216 4988 9280
rect 5052 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5300 9280
rect 4980 8754 5300 9216
rect 4980 8518 5022 8754
rect 5258 8518 5300 8754
rect 4980 8192 5300 8518
rect 4980 8128 4988 8192
rect 5052 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5300 8192
rect 4980 7104 5300 8128
rect 4980 7040 4988 7104
rect 5052 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5300 7104
rect 4980 6170 5300 7040
rect 4980 6016 5022 6170
rect 5258 6016 5300 6170
rect 4980 5952 4988 6016
rect 5292 5952 5300 6016
rect 4980 5934 5022 5952
rect 5258 5934 5300 5952
rect 4980 4928 5300 5934
rect 4980 4864 4988 4928
rect 5052 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5300 4928
rect 4980 3840 5300 4864
rect 4980 3776 4988 3840
rect 5052 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5300 3840
rect 4980 3586 5300 3776
rect 4980 3350 5022 3586
rect 5258 3350 5300 3586
rect 4980 2752 5300 3350
rect 4980 2688 4988 2752
rect 5052 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5300 2752
rect 4980 2128 5300 2688
rect 5640 12000 5960 12560
rect 5640 11936 5648 12000
rect 5712 11998 5728 12000
rect 5792 11998 5808 12000
rect 5872 11998 5888 12000
rect 5952 11936 5960 12000
rect 5640 11762 5682 11936
rect 5918 11762 5960 11936
rect 5640 10912 5960 11762
rect 5640 10848 5648 10912
rect 5712 10848 5728 10912
rect 5792 10848 5808 10912
rect 5872 10848 5888 10912
rect 5952 10848 5960 10912
rect 5640 9824 5960 10848
rect 7671 12544 7991 12560
rect 7671 12480 7679 12544
rect 7743 12480 7759 12544
rect 7823 12480 7839 12544
rect 7903 12480 7919 12544
rect 7983 12480 7991 12544
rect 7671 11456 7991 12480
rect 7671 11392 7679 11456
rect 7743 11392 7759 11456
rect 7823 11392 7839 11456
rect 7903 11392 7919 11456
rect 7983 11392 7991 11456
rect 7671 11338 7991 11392
rect 7671 11102 7713 11338
rect 7949 11102 7991 11338
rect 7671 10368 7991 11102
rect 7671 10304 7679 10368
rect 7743 10304 7759 10368
rect 7823 10304 7839 10368
rect 7903 10304 7919 10368
rect 7983 10304 7991 10368
rect 7419 9892 7485 9893
rect 7419 9828 7420 9892
rect 7484 9828 7485 9892
rect 7419 9827 7485 9828
rect 5640 9760 5648 9824
rect 5712 9760 5728 9824
rect 5792 9760 5808 9824
rect 5872 9760 5888 9824
rect 5952 9760 5960 9824
rect 5640 9414 5960 9760
rect 5640 9178 5682 9414
rect 5918 9178 5960 9414
rect 5640 8736 5960 9178
rect 5640 8672 5648 8736
rect 5712 8672 5728 8736
rect 5792 8672 5808 8736
rect 5872 8672 5888 8736
rect 5952 8672 5960 8736
rect 5640 7648 5960 8672
rect 5640 7584 5648 7648
rect 5712 7584 5728 7648
rect 5792 7584 5808 7648
rect 5872 7584 5888 7648
rect 5952 7584 5960 7648
rect 5640 6830 5960 7584
rect 5640 6594 5682 6830
rect 5918 6594 5960 6830
rect 5640 6560 5960 6594
rect 5640 6496 5648 6560
rect 5712 6496 5728 6560
rect 5792 6496 5808 6560
rect 5872 6496 5888 6560
rect 5952 6496 5960 6560
rect 5640 5472 5960 6496
rect 5640 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5960 5472
rect 5640 4384 5960 5408
rect 5640 4320 5648 4384
rect 5712 4320 5728 4384
rect 5792 4320 5808 4384
rect 5872 4320 5888 4384
rect 5952 4320 5960 4384
rect 5640 4246 5960 4320
rect 5640 4010 5682 4246
rect 5918 4010 5960 4246
rect 5640 3296 5960 4010
rect 5640 3232 5648 3296
rect 5712 3232 5728 3296
rect 5792 3232 5808 3296
rect 5872 3232 5888 3296
rect 5952 3232 5960 3296
rect 5640 2208 5960 3232
rect 7422 2685 7482 9827
rect 7671 9280 7991 10304
rect 7671 9216 7679 9280
rect 7743 9216 7759 9280
rect 7823 9216 7839 9280
rect 7903 9216 7919 9280
rect 7983 9216 7991 9280
rect 7671 8754 7991 9216
rect 7671 8518 7713 8754
rect 7949 8518 7991 8754
rect 7671 8192 7991 8518
rect 7671 8128 7679 8192
rect 7743 8128 7759 8192
rect 7823 8128 7839 8192
rect 7903 8128 7919 8192
rect 7983 8128 7991 8192
rect 7671 7104 7991 8128
rect 7671 7040 7679 7104
rect 7743 7040 7759 7104
rect 7823 7040 7839 7104
rect 7903 7040 7919 7104
rect 7983 7040 7991 7104
rect 7671 6170 7991 7040
rect 7671 6016 7713 6170
rect 7949 6016 7991 6170
rect 7671 5952 7679 6016
rect 7983 5952 7991 6016
rect 7671 5934 7713 5952
rect 7949 5934 7991 5952
rect 7671 4928 7991 5934
rect 7671 4864 7679 4928
rect 7743 4864 7759 4928
rect 7823 4864 7839 4928
rect 7903 4864 7919 4928
rect 7983 4864 7991 4928
rect 7671 3840 7991 4864
rect 7671 3776 7679 3840
rect 7743 3776 7759 3840
rect 7823 3776 7839 3840
rect 7903 3776 7919 3840
rect 7983 3776 7991 3840
rect 7671 3586 7991 3776
rect 7671 3350 7713 3586
rect 7949 3350 7991 3586
rect 7671 2752 7991 3350
rect 7671 2688 7679 2752
rect 7743 2688 7759 2752
rect 7823 2688 7839 2752
rect 7903 2688 7919 2752
rect 7983 2688 7991 2752
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 5640 2144 5648 2208
rect 5712 2144 5728 2208
rect 5792 2144 5808 2208
rect 5872 2144 5888 2208
rect 5952 2144 5960 2208
rect 5640 2128 5960 2144
rect 7671 2128 7991 2688
rect 8331 12000 8651 12560
rect 8331 11936 8339 12000
rect 8403 11998 8419 12000
rect 8483 11998 8499 12000
rect 8563 11998 8579 12000
rect 8643 11936 8651 12000
rect 8331 11762 8373 11936
rect 8609 11762 8651 11936
rect 8331 10912 8651 11762
rect 8331 10848 8339 10912
rect 8403 10848 8419 10912
rect 8483 10848 8499 10912
rect 8563 10848 8579 10912
rect 8643 10848 8651 10912
rect 8331 9824 8651 10848
rect 8331 9760 8339 9824
rect 8403 9760 8419 9824
rect 8483 9760 8499 9824
rect 8563 9760 8579 9824
rect 8643 9760 8651 9824
rect 8331 9414 8651 9760
rect 8331 9178 8373 9414
rect 8609 9178 8651 9414
rect 8331 8736 8651 9178
rect 8331 8672 8339 8736
rect 8403 8672 8419 8736
rect 8483 8672 8499 8736
rect 8563 8672 8579 8736
rect 8643 8672 8651 8736
rect 8331 7648 8651 8672
rect 8331 7584 8339 7648
rect 8403 7584 8419 7648
rect 8483 7584 8499 7648
rect 8563 7584 8579 7648
rect 8643 7584 8651 7648
rect 8331 6830 8651 7584
rect 8331 6594 8373 6830
rect 8609 6594 8651 6830
rect 8331 6560 8651 6594
rect 8331 6496 8339 6560
rect 8403 6496 8419 6560
rect 8483 6496 8499 6560
rect 8563 6496 8579 6560
rect 8643 6496 8651 6560
rect 8331 5472 8651 6496
rect 8331 5408 8339 5472
rect 8403 5408 8419 5472
rect 8483 5408 8499 5472
rect 8563 5408 8579 5472
rect 8643 5408 8651 5472
rect 8331 4384 8651 5408
rect 8331 4320 8339 4384
rect 8403 4320 8419 4384
rect 8483 4320 8499 4384
rect 8563 4320 8579 4384
rect 8643 4320 8651 4384
rect 8331 4246 8651 4320
rect 8331 4010 8373 4246
rect 8609 4010 8651 4246
rect 8331 3296 8651 4010
rect 8331 3232 8339 3296
rect 8403 3232 8419 3296
rect 8483 3232 8499 3296
rect 8563 3232 8579 3296
rect 8643 3232 8651 3296
rect 8331 2208 8651 3232
rect 8331 2144 8339 2208
rect 8403 2144 8419 2208
rect 8483 2144 8499 2208
rect 8563 2144 8579 2208
rect 8643 2144 8651 2208
rect 8331 2128 8651 2144
rect 10362 12544 10682 12560
rect 10362 12480 10370 12544
rect 10434 12480 10450 12544
rect 10514 12480 10530 12544
rect 10594 12480 10610 12544
rect 10674 12480 10682 12544
rect 10362 11456 10682 12480
rect 10362 11392 10370 11456
rect 10434 11392 10450 11456
rect 10514 11392 10530 11456
rect 10594 11392 10610 11456
rect 10674 11392 10682 11456
rect 10362 11338 10682 11392
rect 10362 11102 10404 11338
rect 10640 11102 10682 11338
rect 10362 10368 10682 11102
rect 10362 10304 10370 10368
rect 10434 10304 10450 10368
rect 10514 10304 10530 10368
rect 10594 10304 10610 10368
rect 10674 10304 10682 10368
rect 10362 9280 10682 10304
rect 10362 9216 10370 9280
rect 10434 9216 10450 9280
rect 10514 9216 10530 9280
rect 10594 9216 10610 9280
rect 10674 9216 10682 9280
rect 10362 8754 10682 9216
rect 10362 8518 10404 8754
rect 10640 8518 10682 8754
rect 10362 8192 10682 8518
rect 10362 8128 10370 8192
rect 10434 8128 10450 8192
rect 10514 8128 10530 8192
rect 10594 8128 10610 8192
rect 10674 8128 10682 8192
rect 10362 7104 10682 8128
rect 10362 7040 10370 7104
rect 10434 7040 10450 7104
rect 10514 7040 10530 7104
rect 10594 7040 10610 7104
rect 10674 7040 10682 7104
rect 10362 6170 10682 7040
rect 10362 6016 10404 6170
rect 10640 6016 10682 6170
rect 10362 5952 10370 6016
rect 10674 5952 10682 6016
rect 10362 5934 10404 5952
rect 10640 5934 10682 5952
rect 10362 4928 10682 5934
rect 10362 4864 10370 4928
rect 10434 4864 10450 4928
rect 10514 4864 10530 4928
rect 10594 4864 10610 4928
rect 10674 4864 10682 4928
rect 10362 3840 10682 4864
rect 10362 3776 10370 3840
rect 10434 3776 10450 3840
rect 10514 3776 10530 3840
rect 10594 3776 10610 3840
rect 10674 3776 10682 3840
rect 10362 3586 10682 3776
rect 10362 3350 10404 3586
rect 10640 3350 10682 3586
rect 10362 2752 10682 3350
rect 10362 2688 10370 2752
rect 10434 2688 10450 2752
rect 10514 2688 10530 2752
rect 10594 2688 10610 2752
rect 10674 2688 10682 2752
rect 10362 2128 10682 2688
rect 11022 12000 11342 12560
rect 11022 11936 11030 12000
rect 11094 11998 11110 12000
rect 11174 11998 11190 12000
rect 11254 11998 11270 12000
rect 11334 11936 11342 12000
rect 11022 11762 11064 11936
rect 11300 11762 11342 11936
rect 11022 10912 11342 11762
rect 11022 10848 11030 10912
rect 11094 10848 11110 10912
rect 11174 10848 11190 10912
rect 11254 10848 11270 10912
rect 11334 10848 11342 10912
rect 11022 9824 11342 10848
rect 11022 9760 11030 9824
rect 11094 9760 11110 9824
rect 11174 9760 11190 9824
rect 11254 9760 11270 9824
rect 11334 9760 11342 9824
rect 11022 9414 11342 9760
rect 11022 9178 11064 9414
rect 11300 9178 11342 9414
rect 11022 8736 11342 9178
rect 11022 8672 11030 8736
rect 11094 8672 11110 8736
rect 11174 8672 11190 8736
rect 11254 8672 11270 8736
rect 11334 8672 11342 8736
rect 11022 7648 11342 8672
rect 11022 7584 11030 7648
rect 11094 7584 11110 7648
rect 11174 7584 11190 7648
rect 11254 7584 11270 7648
rect 11334 7584 11342 7648
rect 11022 6830 11342 7584
rect 11022 6594 11064 6830
rect 11300 6594 11342 6830
rect 11022 6560 11342 6594
rect 11022 6496 11030 6560
rect 11094 6496 11110 6560
rect 11174 6496 11190 6560
rect 11254 6496 11270 6560
rect 11334 6496 11342 6560
rect 11022 5472 11342 6496
rect 11022 5408 11030 5472
rect 11094 5408 11110 5472
rect 11174 5408 11190 5472
rect 11254 5408 11270 5472
rect 11334 5408 11342 5472
rect 11022 4384 11342 5408
rect 11022 4320 11030 4384
rect 11094 4320 11110 4384
rect 11174 4320 11190 4384
rect 11254 4320 11270 4384
rect 11334 4320 11342 4384
rect 11022 4246 11342 4320
rect 11022 4010 11064 4246
rect 11300 4010 11342 4246
rect 11022 3296 11342 4010
rect 11022 3232 11030 3296
rect 11094 3232 11110 3296
rect 11174 3232 11190 3296
rect 11254 3232 11270 3296
rect 11334 3232 11342 3296
rect 11022 2208 11342 3232
rect 11022 2144 11030 2208
rect 11094 2144 11110 2208
rect 11174 2144 11190 2208
rect 11254 2144 11270 2208
rect 11334 2144 11342 2208
rect 11022 2128 11342 2144
<< via4 >>
rect 2331 11102 2567 11338
rect 2331 8518 2567 8754
rect 2331 6016 2567 6170
rect 2331 5952 2361 6016
rect 2361 5952 2377 6016
rect 2377 5952 2441 6016
rect 2441 5952 2457 6016
rect 2457 5952 2521 6016
rect 2521 5952 2537 6016
rect 2537 5952 2567 6016
rect 2331 5934 2567 5952
rect 2331 3350 2567 3586
rect 2991 11936 3021 11998
rect 3021 11936 3037 11998
rect 3037 11936 3101 11998
rect 3101 11936 3117 11998
rect 3117 11936 3181 11998
rect 3181 11936 3197 11998
rect 3197 11936 3227 11998
rect 2991 11762 3227 11936
rect 2991 9178 3227 9414
rect 2991 6594 3227 6830
rect 2991 4010 3227 4246
rect 5022 11102 5258 11338
rect 5022 8518 5258 8754
rect 5022 6016 5258 6170
rect 5022 5952 5052 6016
rect 5052 5952 5068 6016
rect 5068 5952 5132 6016
rect 5132 5952 5148 6016
rect 5148 5952 5212 6016
rect 5212 5952 5228 6016
rect 5228 5952 5258 6016
rect 5022 5934 5258 5952
rect 5022 3350 5258 3586
rect 5682 11936 5712 11998
rect 5712 11936 5728 11998
rect 5728 11936 5792 11998
rect 5792 11936 5808 11998
rect 5808 11936 5872 11998
rect 5872 11936 5888 11998
rect 5888 11936 5918 11998
rect 5682 11762 5918 11936
rect 7713 11102 7949 11338
rect 5682 9178 5918 9414
rect 5682 6594 5918 6830
rect 5682 4010 5918 4246
rect 7713 8518 7949 8754
rect 7713 6016 7949 6170
rect 7713 5952 7743 6016
rect 7743 5952 7759 6016
rect 7759 5952 7823 6016
rect 7823 5952 7839 6016
rect 7839 5952 7903 6016
rect 7903 5952 7919 6016
rect 7919 5952 7949 6016
rect 7713 5934 7949 5952
rect 7713 3350 7949 3586
rect 8373 11936 8403 11998
rect 8403 11936 8419 11998
rect 8419 11936 8483 11998
rect 8483 11936 8499 11998
rect 8499 11936 8563 11998
rect 8563 11936 8579 11998
rect 8579 11936 8609 11998
rect 8373 11762 8609 11936
rect 8373 9178 8609 9414
rect 8373 6594 8609 6830
rect 8373 4010 8609 4246
rect 10404 11102 10640 11338
rect 10404 8518 10640 8754
rect 10404 6016 10640 6170
rect 10404 5952 10434 6016
rect 10434 5952 10450 6016
rect 10450 5952 10514 6016
rect 10514 5952 10530 6016
rect 10530 5952 10594 6016
rect 10594 5952 10610 6016
rect 10610 5952 10640 6016
rect 10404 5934 10640 5952
rect 10404 3350 10640 3586
rect 11064 11936 11094 11998
rect 11094 11936 11110 11998
rect 11110 11936 11174 11998
rect 11174 11936 11190 11998
rect 11190 11936 11254 11998
rect 11254 11936 11270 11998
rect 11270 11936 11300 11998
rect 11064 11762 11300 11936
rect 11064 9178 11300 9414
rect 11064 6594 11300 6830
rect 11064 4010 11300 4246
<< metal5 >>
rect 1056 11998 11916 12040
rect 1056 11762 2991 11998
rect 3227 11762 5682 11998
rect 5918 11762 8373 11998
rect 8609 11762 11064 11998
rect 11300 11762 11916 11998
rect 1056 11720 11916 11762
rect 1056 11338 11916 11380
rect 1056 11102 2331 11338
rect 2567 11102 5022 11338
rect 5258 11102 7713 11338
rect 7949 11102 10404 11338
rect 10640 11102 11916 11338
rect 1056 11060 11916 11102
rect 1056 9414 11916 9456
rect 1056 9178 2991 9414
rect 3227 9178 5682 9414
rect 5918 9178 8373 9414
rect 8609 9178 11064 9414
rect 11300 9178 11916 9414
rect 1056 9136 11916 9178
rect 1056 8754 11916 8796
rect 1056 8518 2331 8754
rect 2567 8518 5022 8754
rect 5258 8518 7713 8754
rect 7949 8518 10404 8754
rect 10640 8518 11916 8754
rect 1056 8476 11916 8518
rect 1056 6830 11916 6872
rect 1056 6594 2991 6830
rect 3227 6594 5682 6830
rect 5918 6594 8373 6830
rect 8609 6594 11064 6830
rect 11300 6594 11916 6830
rect 1056 6552 11916 6594
rect 1056 6170 11916 6212
rect 1056 5934 2331 6170
rect 2567 5934 5022 6170
rect 5258 5934 7713 6170
rect 7949 5934 10404 6170
rect 10640 5934 11916 6170
rect 1056 5892 11916 5934
rect 1056 4246 11916 4288
rect 1056 4010 2991 4246
rect 3227 4010 5682 4246
rect 5918 4010 8373 4246
rect 8609 4010 11064 4246
rect 11300 4010 11916 4246
rect 1056 3968 11916 4010
rect 1056 3586 11916 3628
rect 1056 3350 2331 3586
rect 2567 3350 5022 3586
rect 5258 3350 7713 3586
rect 7949 3350 10404 3586
rect 10640 3350 11916 3586
rect 1056 3308 11916 3350
use sky130_fd_sc_hd__inv_2  _151_
timestamp 0
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 0
transform -1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 0
transform -1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 0
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 0
transform -1 0 6164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 0
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 0
transform -1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _159_
timestamp 0
transform 1 0 5060 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 0
transform -1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 0
transform 1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _162_
timestamp 0
transform 1 0 4140 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _163_
timestamp 0
transform -1 0 4876 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _164_
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _165_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_4  _166_
timestamp 0
transform 1 0 5060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _167_
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _168_
timestamp 0
transform 1 0 10212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _169_
timestamp 0
transform 1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _170_
timestamp 0
transform -1 0 11316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _171_
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _172_
timestamp 0
transform -1 0 10856 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _173_
timestamp 0
transform -1 0 9200 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _174_
timestamp 0
transform 1 0 7268 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _175_
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _176_
timestamp 0
transform -1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _177_
timestamp 0
transform 1 0 9476 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _178_
timestamp 0
transform -1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _179_
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _180_
timestamp 0
transform -1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 0
transform -1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _182_
timestamp 0
transform 1 0 7820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _183_
timestamp 0
transform 1 0 7268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _184_
timestamp 0
transform -1 0 8280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _185_
timestamp 0
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_4  _186_
timestamp 0
transform 1 0 6808 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__o21a_1  _187_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _188_
timestamp 0
transform -1 0 4692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _189_
timestamp 0
transform -1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _190_
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _191_
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _192_
timestamp 0
transform -1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 0
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 0
transform -1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 0
transform -1 0 10764 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 0
transform -1 0 3312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _197_
timestamp 0
transform -1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _198_
timestamp 0
transform -1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _199_
timestamp 0
transform -1 0 2852 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 0
transform -1 0 3312 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 0
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _203_
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _204_
timestamp 0
transform 1 0 1748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _205_
timestamp 0
transform 1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _206_
timestamp 0
transform 1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _207_
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _208_
timestamp 0
transform 1 0 2024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _209_
timestamp 0
transform 1 0 2208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_4  _210_
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_1  _211_
timestamp 0
transform 1 0 1932 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 0
transform 1 0 3312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _213_
timestamp 0
transform -1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _214_
timestamp 0
transform 1 0 2760 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _215_
timestamp 0
transform 1 0 5336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _216_
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 0
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _219_
timestamp 0
transform -1 0 6992 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _220_
timestamp 0
transform -1 0 10856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _221_
timestamp 0
transform -1 0 11316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _222_
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 0
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _224_
timestamp 0
transform 1 0 9936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _225_
timestamp 0
transform -1 0 11500 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _226_
timestamp 0
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 0
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _229_
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _230_
timestamp 0
transform -1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _231_
timestamp 0
transform -1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _232_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _233_
timestamp 0
transform -1 0 8556 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _234_
timestamp 0
transform -1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _235_
timestamp 0
transform 1 0 5520 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 0
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 0
transform 1 0 4324 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _238_
timestamp 0
transform -1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _239_
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _240_
timestamp 0
transform -1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _241_
timestamp 0
transform 1 0 4784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 0
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _243_
timestamp 0
transform 1 0 9844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _244_
timestamp 0
transform 1 0 10120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _245_
timestamp 0
transform 1 0 9752 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _246_
timestamp 0
transform 1 0 10304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _248_
timestamp 0
transform -1 0 11040 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _250_
timestamp 0
transform 1 0 10488 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _251_
timestamp 0
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _252_
timestamp 0
transform -1 0 7912 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _253_
timestamp 0
transform -1 0 6256 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _254_
timestamp 0
transform 1 0 7176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _255_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_4  _256_
timestamp 0
transform -1 0 8096 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_2  _257_
timestamp 0
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _258_
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _259_
timestamp 0
transform 1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 0
transform 1 0 6992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _261_
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _262_
timestamp 0
transform 1 0 7452 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _263_
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _264_
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _265_
timestamp 0
transform 1 0 3864 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _266_
timestamp 0
transform -1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _267_
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _268_
timestamp 0
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _269_
timestamp 0
transform 1 0 5152 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _270_
timestamp 0
transform -1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _271_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _272_
timestamp 0
transform -1 0 5980 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _273_
timestamp 0
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _274_
timestamp 0
transform -1 0 6164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _275_
timestamp 0
transform -1 0 10212 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _276_
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _277_
timestamp 0
transform 1 0 9016 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _278_
timestamp 0
transform 1 0 9292 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 0
transform -1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _280_
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _281_
timestamp 0
transform -1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _282_
timestamp 0
transform -1 0 9844 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 0
transform -1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _284_
timestamp 0
transform 1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _285_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _286_
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _287_
timestamp 0
transform -1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _288_
timestamp 0
transform 1 0 7452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _289_
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _290_
timestamp 0
transform 1 0 3312 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _291_
timestamp 0
transform -1 0 8096 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _292_
timestamp 0
transform 1 0 6808 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _293_
timestamp 0
transform 1 0 7636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _294_
timestamp 0
transform -1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _295_
timestamp 0
transform -1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _296_
timestamp 0
transform -1 0 9108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _297_
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _298_
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _299_
timestamp 0
transform -1 0 8372 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 0
transform -1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 0
transform -1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _302_
timestamp 0
transform 1 0 1564 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _303_
timestamp 0
transform -1 0 5888 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _304_
timestamp 0
transform 1 0 2392 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _305_
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _306_
timestamp 0
transform -1 0 4508 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _307_
timestamp 0
transform -1 0 3680 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _308_
timestamp 0
transform -1 0 3496 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _309_
timestamp 0
transform -1 0 3496 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform -1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 0
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_71
timestamp 0
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_93
timestamp 0
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_104
timestamp 0
transform 1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_64
timestamp 0
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_86
timestamp 0
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_90
timestamp 0
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_97
timestamp 0
transform 1 0 10028 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_108
timestamp 0
transform 1 0 11040 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_91
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_102
timestamp 0
transform 1 0 10488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_9
timestamp 0
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_13
timestamp 0
transform 1 0 2300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_40
timestamp 0
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_87
timestamp 0
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_57
timestamp 0
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_69
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 0
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_93
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_113
timestamp 0
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_9
timestamp 0
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_13
timestamp 0
transform 1 0 2300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_37
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_45
timestamp 0
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_84
timestamp 0
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_96
timestamp 0
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_100
timestamp 0
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_104
timestamp 0
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_108
timestamp 0
transform 1 0 11040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 0
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_93
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_99
timestamp 0
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_108
timestamp 0
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_63
timestamp 0
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_84
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_88
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_96
timestamp 0
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 0
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_34
timestamp 0
transform 1 0 4232 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_55
timestamp 0
transform 1 0 6164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_67
timestamp 0
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_91
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_95
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_100
timestamp 0
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_112
timestamp 0
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_24
timestamp 0
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_32
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_65
timestamp 0
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_74
timestamp 0
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_86
timestamp 0
transform 1 0 9016 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_98
timestamp 0
transform 1 0 10120 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_38
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_46
timestamp 0
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_12
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_31
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_64
timestamp 0
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_72
timestamp 0
transform 1 0 7728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_84
timestamp 0
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 0
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_51
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_63
timestamp 0
transform 1 0 6900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_71
timestamp 0
transform 1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 0
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_91
timestamp 0
transform 1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_108
timestamp 0
transform 1 0 11040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_16
timestamp 0
transform 1 0 2576 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_29
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_33
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_41
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_47
timestamp 0
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_63
timestamp 0
transform 1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_87
timestamp 0
transform 1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_95
timestamp 0
transform 1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 0
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_6
timestamp 0
transform 1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_40
timestamp 0
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_50
timestamp 0
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_62
timestamp 0
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 0
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_103
timestamp 0
transform 1 0 10580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_6
timestamp 0
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_24
timestamp 0
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_36
timestamp 0
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_48
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_16
timestamp 0
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_38
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_55
timestamp 0
transform 1 0 6164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_61
timestamp 0
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 0
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_6
timestamp 0
transform 1 0 1656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_13
timestamp 0
transform 1 0 2300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_47
timestamp 0
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_88
timestamp 0
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_16
timestamp 0
transform 1 0 2576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_20
timestamp 0
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_37
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_51
timestamp 0
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_55
timestamp 0
transform 1 0 6164 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_57
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_62
timestamp 0
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 0
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_75
timestamp 0
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_90
timestamp 0
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_94
timestamp 0
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_105
timestamp 0
transform 1 0 10764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_111
timestamp 0
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_113
timestamp 0
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform -1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 0
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 0
transform -1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform -1 0 11592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 0
transform -1 0 11408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform -1 0 8740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 0
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 0
transform 1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 0
transform 1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 0
transform -1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 0
transform -1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 0
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 0
transform -1 0 11408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 0
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 0
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 0
transform -1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 0
transform -1 0 11408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 0
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 0
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 0
transform 1 0 9844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 0
transform -1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 0
transform -1 0 5796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 0
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 0
transform -1 0 1932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 11868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 11868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 1 11968
box -38 -48 130 592
<< labels >>
rlabel metal1 s 6486 11968 6486 11968 4 VGND
rlabel metal1 s 6486 12512 6486 12512 4 VPWR
rlabel metal2 s 4646 3876 4646 3876 4 _000_
rlabel metal1 s 4876 3162 4876 3162 4 _001_
rlabel metal1 s 5428 4114 5428 4114 4 _002_
rlabel metal1 s 5658 4250 5658 4250 4 _003_
rlabel metal1 s 4469 3094 4469 3094 4 _004_
rlabel metal1 s 3089 3434 3089 3434 4 _005_
rlabel metal1 s 2905 2346 2905 2346 4 _006_
rlabel metal1 s 2744 5610 2744 5610 4 _007_
rlabel metal2 s 7682 4522 7682 4522 4 _008_
rlabel metal1 s 6081 3706 6081 3706 4 _009_
rlabel metal2 s 2162 5168 2162 5168 4 _010_
rlabel metal1 s 2346 5236 2346 5236 4 _011_
rlabel metal2 s 4186 3978 4186 3978 4 _012_
rlabel metal2 s 3358 4063 3358 4063 4 _013_
rlabel metal1 s 3312 2346 3312 2346 4 _014_
rlabel metal1 s 4646 5610 4646 5610 4 _015_
rlabel metal1 s 2300 7310 2300 7310 4 _016_
rlabel metal1 s 2852 7514 2852 7514 4 _017_
rlabel metal3 s 3266 7973 3266 7973 4 _018_
rlabel metal1 s 3634 7718 3634 7718 4 _019_
rlabel metal1 s 2622 8534 2622 8534 4 _020_
rlabel metal1 s 2208 9010 2208 9010 4 _021_
rlabel metal1 s 2622 8398 2622 8398 4 _022_
rlabel metal1 s 2116 10030 2116 10030 4 _023_
rlabel metal1 s 2162 7514 2162 7514 4 _024_
rlabel metal1 s 2668 8058 2668 8058 4 _025_
rlabel metal2 s 3358 9554 3358 9554 4 _026_
rlabel metal2 s 9614 7514 9614 7514 4 _027_
rlabel metal2 s 2806 10982 2806 10982 4 _028_
rlabel metal1 s 3680 11186 3680 11186 4 _029_
rlabel metal1 s 3404 10778 3404 10778 4 _030_
rlabel metal1 s 3128 9554 3128 9554 4 _031_
rlabel metal1 s 9200 7854 9200 7854 4 _032_
rlabel metal1 s 5842 6800 5842 6800 4 _033_
rlabel metal1 s 7084 2890 7084 2890 4 _034_
rlabel metal1 s 5934 2992 5934 2992 4 _035_
rlabel metal1 s 7452 3094 7452 3094 4 _036_
rlabel metal2 s 10166 3978 10166 3978 4 _037_
rlabel metal1 s 10304 4114 10304 4114 4 _038_
rlabel metal1 s 10028 3162 10028 3162 4 _039_
rlabel metal1 s 9982 4080 9982 4080 4 _040_
rlabel metal2 s 10258 3808 10258 3808 4 _041_
rlabel metal1 s 10580 3570 10580 3570 4 _042_
rlabel metal1 s 8141 3026 8141 3026 4 _043_
rlabel metal1 s 7498 3604 7498 3604 4 _044_
rlabel metal2 s 7314 3570 7314 3570 4 _045_
rlabel metal2 s 8234 3230 8234 3230 4 _046_
rlabel metal1 s 8004 2822 8004 2822 4 _047_
rlabel metal2 s 7498 3196 7498 3196 4 _048_
rlabel metal1 s 8510 3604 8510 3604 4 _049_
rlabel metal2 s 8323 6290 8323 6290 4 _050_
rlabel metal1 s 6072 6154 6072 6154 4 _051_
rlabel metal1 s 4462 6426 4462 6426 4 _052_
rlabel metal1 s 5106 6732 5106 6732 4 _053_
rlabel metal1 s 5290 6902 5290 6902 4 _054_
rlabel metal1 s 5290 6800 5290 6800 4 _055_
rlabel metal2 s 8740 5202 8740 5202 4 _056_
rlabel metal2 s 5290 6460 5290 6460 4 _057_
rlabel metal1 s 2369 10098 2369 10098 4 _058_
rlabel metal1 s 10488 8602 10488 8602 4 _059_
rlabel metal1 s 10608 8942 10608 8942 4 _060_
rlabel metal1 s 10304 8942 10304 8942 4 _061_
rlabel metal1 s 11086 8602 11086 8602 4 _062_
rlabel metal1 s 10812 6290 10812 6290 4 _063_
rlabel metal1 s 11178 8466 11178 8466 4 _064_
rlabel metal1 s 10902 6800 10902 6800 4 _065_
rlabel metal1 s 11270 6970 11270 6970 4 _066_
rlabel metal1 s 9384 8398 9384 8398 4 _067_
rlabel metal1 s 7452 7514 7452 7514 4 _068_
rlabel metal1 s 7406 8432 7406 8432 4 _069_
rlabel metal1 s 7176 7922 7176 7922 4 _070_
rlabel metal2 s 6946 8058 6946 8058 4 _071_
rlabel metal1 s 7636 6358 7636 6358 4 _072_
rlabel metal1 s 8050 6358 8050 6358 4 _073_
rlabel metal1 s 6946 2822 6946 2822 4 _074_
rlabel metal1 s 5796 5882 5796 5882 4 _075_
rlabel metal1 s 7751 5202 7751 5202 4 _076_
rlabel metal2 s 8234 5746 8234 5746 4 _077_
rlabel metal2 s 5290 8636 5290 8636 4 _078_
rlabel metal2 s 6118 8194 6118 8194 4 _079_
rlabel metal1 s 4462 8058 4462 8058 4 _080_
rlabel metal1 s 5801 4590 5801 4590 4 _081_
rlabel metal1 s 5428 3162 5428 3162 4 _082_
rlabel metal1 s 5612 5814 5612 5814 4 _083_
rlabel metal1 s 5566 5712 5566 5712 4 _084_
rlabel metal1 s 4830 5678 4830 5678 4 _085_
rlabel metal2 s 6025 5202 6025 5202 4 _086_
rlabel metal1 s 6072 3162 6072 3162 4 _087_
rlabel metal1 s 9660 5882 9660 5882 4 _088_
rlabel metal1 s 10258 6154 10258 6154 4 _089_
rlabel metal2 s 9798 6460 9798 6460 4 _090_
rlabel metal1 s 8417 5202 8417 5202 4 _091_
rlabel metal2 s 10074 4998 10074 4998 4 _092_
rlabel metal1 s 8510 5168 8510 5168 4 _093_
rlabel metal2 s 9246 8160 9246 8160 4 _094_
rlabel metal2 s 9338 8126 9338 8126 4 _095_
rlabel metal1 s 9430 7820 9430 7820 4 _096_
rlabel metal2 s 8693 6290 8693 6290 4 _097_
rlabel metal1 s 8786 6256 8786 6256 4 _098_
rlabel metal1 s 7820 9418 7820 9418 4 _099_
rlabel metal1 s 7912 9486 7912 9486 4 _100_
rlabel metal1 s 7590 9486 7590 9486 4 _101_
rlabel metal2 s 7848 4590 7848 4590 4 _102_
rlabel metal1 s 7544 4590 7544 4590 4 _103_
rlabel metal1 s 8188 9078 8188 9078 4 _104_
rlabel metal1 s 8878 9010 8878 9010 4 _105_
rlabel metal1 s 8556 8942 8556 8942 4 _106_
rlabel metal2 s 8160 4114 8160 4114 4 _107_
rlabel metal1 s 8510 4114 8510 4114 4 _108_
rlabel metal1 s 6486 3366 6486 3366 4 _109_
rlabel metal1 s 5658 8432 5658 8432 4 _110_
rlabel metal1 s 5658 11186 5658 11186 4 _111_
rlabel metal2 s 5934 8415 5934 8415 4 _112_
rlabel metal1 s 10764 4998 10764 4998 4 _113_
rlabel metal1 s 4738 11050 4738 11050 4 _114_
rlabel metal2 s 4738 10370 4738 10370 4 _115_
rlabel metal1 s 6302 11730 6302 11730 4 _116_
rlabel metal1 s 5842 11118 5842 11118 4 _117_
rlabel metal1 s 6164 10642 6164 10642 4 _118_
rlabel metal1 s 10534 11084 10534 11084 4 _119_
rlabel metal2 s 10902 11220 10902 11220 4 _120_
rlabel metal1 s 10074 11152 10074 11152 4 _121_
rlabel metal2 s 10626 11186 10626 11186 4 _122_
rlabel metal1 s 10488 10778 10488 10778 4 _123_
rlabel metal1 s 9706 11152 9706 11152 4 _124_
rlabel metal2 s 8234 11900 8234 11900 4 _125_
rlabel metal2 s 8050 12002 8050 12002 4 _126_
rlabel metal2 s 7958 11900 7958 11900 4 _127_
rlabel metal2 s 9798 11730 9798 11730 4 _128_
rlabel metal1 s 6762 10506 6762 10506 4 _129_
rlabel metal1 s 5428 10710 5428 10710 4 _130_
rlabel metal1 s 6716 10030 6716 10030 4 _131_
rlabel metal2 s 10074 6528 10074 6528 4 _132_
rlabel metal2 s 7958 10948 7958 10948 4 _133_
rlabel metal2 s 7130 11356 7130 11356 4 _134_
rlabel metal1 s 7804 10710 7804 10710 4 _135_
rlabel metal2 s 9614 6188 9614 6188 4 _136_
rlabel metal1 s 6900 9554 6900 9554 4 _137_
rlabel metal1 s 6992 9486 6992 9486 4 _138_
rlabel metal1 s 6118 9520 6118 9520 4 _139_
rlabel metal2 s 3542 11356 3542 11356 4 _140_
rlabel metal1 s 2530 11322 2530 11322 4 _141_
rlabel metal1 s 2116 10982 2116 10982 4 _142_
rlabel metal2 s 1978 11390 1978 11390 4 _143_
rlabel metal2 s 2898 10948 2898 10948 4 _144_
rlabel metal1 s 11040 5882 11040 5882 4 _145_
rlabel metal2 s 10810 4386 10810 4386 4 _146_
rlabel metal1 s 3818 11118 3818 11118 4 _147_
rlabel metal1 s 3220 10030 3220 10030 4 _148_
rlabel metal1 s 3358 11084 3358 11084 4 _149_
rlabel metal1 s 1932 7786 1932 7786 4 _150_
rlabel metal3 s 1004 4148 1004 4148 4 clk
rlabel metal1 s 4370 2414 4370 2414 4 clknet_0_clk
rlabel metal1 s 3542 2482 3542 2482 4 clknet_1_0__leaf_clk
rlabel metal2 s 2714 5984 2714 5984 4 clknet_1_1__leaf_clk
rlabel metal2 s 10350 1027 10350 1027 4 input_data_0[0]
rlabel metal2 s 6539 14484 6539 14484 4 input_data_0[1]
rlabel metal3 s 820 10948 820 10948 4 input_data_0[2]
rlabel metal2 s 12926 1554 12926 1554 4 input_data_0[3]
rlabel metal1 s 10350 2448 10350 2448 4 input_data_0[4]
rlabel metal2 s 11546 9809 11546 9809 4 input_data_0[5]
rlabel metal1 s 2346 12240 2346 12240 4 input_data_0[6]
rlabel metal3 s 866 12308 866 12308 4 input_data_0[7]
rlabel metal2 s 10304 12716 10304 12716 4 input_data_1[0]
rlabel metal2 s 7774 1588 7774 1588 4 input_data_1[1]
rlabel metal2 s 11546 11033 11546 11033 4 input_data_1[2]
rlabel metal2 s 11362 2907 11362 2907 4 input_data_1[3]
rlabel metal2 s 2622 1435 2622 1435 4 input_data_1[4]
rlabel metal3 s 1050 9588 1050 9588 4 input_data_1[5]
rlabel metal3 s 1050 6868 1050 6868 4 input_data_1[6]
rlabel metal2 s 8694 12410 8694 12410 4 input_data_1[7]
rlabel metal1 s 11224 11866 11224 11866 4 input_data_2[0]
rlabel metal3 s 1050 8228 1050 8228 4 input_data_2[1]
rlabel metal1 s 10534 11696 10534 11696 4 input_data_2[2]
rlabel metal2 s 2714 12801 2714 12801 4 input_data_2[3]
rlabel metal2 s 46 1860 46 1860 4 input_data_2[4]
rlabel metal3 s 820 2788 820 2788 4 input_data_2[5]
rlabel metal2 s 11546 8041 11546 8041 4 input_data_2[6]
rlabel metal1 s 1380 11730 1380 11730 4 input_data_2[7]
rlabel metal3 s 1050 1428 1050 1428 4 input_data_3[0]
rlabel metal2 s 11638 1588 11638 1588 4 input_data_3[1]
rlabel metal1 s 9108 12206 9108 12206 4 input_data_3[2]
rlabel metal1 s 11408 5202 11408 5202 4 input_data_3[3]
rlabel metal2 s 1334 1894 1334 1894 4 input_data_3[4]
rlabel metal2 s 3910 1163 3910 1163 4 input_data_3[5]
rlabel metal2 s 5198 1588 5198 1588 4 input_data_3[6]
rlabel metal2 s 11546 5593 11546 5593 4 input_data_3[7]
rlabel metal1 s 10212 2618 10212 2618 4 net1
rlabel metal1 s 7682 2618 7682 2618 4 net10
rlabel metal1 s 10304 10166 10304 10166 4 net11
rlabel metal1 s 10902 5610 10902 5610 4 net12
rlabel metal2 s 4370 10081 4370 10081 4 net13
rlabel metal1 s 4554 9962 4554 9962 4 net14
rlabel metal2 s 1610 7038 1610 7038 4 net15
rlabel metal2 s 5566 12104 5566 12104 4 net16
rlabel metal3 s 4278 11067 4278 11067 4 net17
rlabel metal2 s 1702 9962 1702 9962 4 net18
rlabel metal2 s 9706 9894 9706 9894 4 net19
rlabel metal2 s 8326 9350 8326 9350 4 net2
rlabel metal1 s 9292 6766 9292 6766 4 net20
rlabel metal1 s 1748 7854 1748 7854 4 net21
rlabel metal1 s 1840 7310 1840 7310 4 net22
rlabel metal1 s 3634 7888 3634 7888 4 net23
rlabel metal1 s 1748 9350 1748 9350 4 net24
rlabel metal3 s 1610 3995 1610 3995 4 net25
rlabel metal1 s 11316 2618 11316 2618 4 net26
rlabel metal1 s 8786 6358 8786 6358 4 net27
rlabel metal2 s 11270 4794 11270 4794 4 net28
rlabel metal2 s 2622 3111 2622 3111 4 net29
rlabel metal2 s 1886 10234 1886 10234 4 net3
rlabel metal3 s 2346 2907 2346 2907 4 net30
rlabel metal1 s 7314 2414 7314 2414 4 net31
rlabel metal1 s 8878 3502 8878 3502 4 net32
rlabel metal1 s 6164 4114 6164 4114 4 net33
rlabel metal2 s 6946 2587 6946 2587 4 net34
rlabel metal1 s 10028 9078 10028 9078 4 net35
rlabel metal1 s 7314 6154 7314 6154 4 net36
rlabel metal1 s 4324 12206 4324 12206 4 net37
rlabel metal1 s 5980 12138 5980 12138 4 net38
rlabel metal1 s 7912 3026 7912 3026 4 net39
rlabel metal1 s 10856 2618 10856 2618 4 net4
rlabel metal2 s 7130 3553 7130 3553 4 net40
rlabel metal1 s 4462 11764 4462 11764 4 net41
rlabel metal1 s 10856 2550 10856 2550 4 net5
rlabel metal1 s 7084 7378 7084 7378 4 net6
rlabel metal1 s 3726 12342 3726 12342 4 net7
rlabel metal2 s 6578 10812 6578 10812 4 net8
rlabel metal1 s 9246 11526 9246 11526 4 net9
rlabel metal2 s 6486 1554 6486 1554 4 output_data[0]
rlabel metal3 s 11922 13668 11922 13668 4 output_data[1]
rlabel metal1 s 11592 12410 11592 12410 4 output_data[2]
rlabel metal1 s 4002 12410 4002 12410 4 output_data[3]
rlabel metal2 s 5290 13260 5290 13260 4 output_data[4]
rlabel metal2 s 9062 1520 9062 1520 4 output_data[5]
rlabel metal3 s 820 5508 820 5508 4 output_data[6]
rlabel metal3 s 1096 13668 1096 13668 4 output_data[7]
rlabel metal2 s 11270 7123 11270 7123 4 reset
flabel metal5 s 1056 11720 11916 12040 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 9136 11916 9456 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6552 11916 6872 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3968 11916 4288 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 11022 2128 11342 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8331 2128 8651 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5640 2128 5960 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2949 2128 3269 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 11060 11916 11380 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8476 11916 8796 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5892 11916 6212 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3308 11916 3628 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 10362 2128 10682 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7671 2128 7991 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4980 2128 5300 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2289 2128 2609 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 4088 800 4208 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 input_data_0[0]
port 4 nsew
flabel metal2 s 6458 14397 6514 15197 0 FreeSans 280 90 0 0 input_data_0[1]
port 5 nsew
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 input_data_0[2]
port 6 nsew
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 input_data_0[3]
port 7 nsew
flabel metal3 s 12253 1368 13053 1488 0 FreeSans 600 0 0 0 input_data_0[4]
port 8 nsew
flabel metal3 s 12253 9528 13053 9648 0 FreeSans 600 0 0 0 input_data_0[5]
port 9 nsew
flabel metal2 s 18 14397 74 15197 0 FreeSans 280 90 0 0 input_data_0[6]
port 10 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 input_data_0[7]
port 11 nsew
flabel metal2 s 10322 14397 10378 15197 0 FreeSans 280 90 0 0 input_data_1[0]
port 12 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 input_data_1[1]
port 13 nsew
flabel metal3 s 12253 10888 13053 11008 0 FreeSans 600 0 0 0 input_data_1[2]
port 14 nsew
flabel metal3 s 12253 2728 13053 2848 0 FreeSans 600 0 0 0 input_data_1[3]
port 15 nsew
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 input_data_1[4]
port 16 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 input_data_1[5]
port 17 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 input_data_1[6]
port 18 nsew
flabel metal2 s 7746 14397 7802 15197 0 FreeSans 280 90 0 0 input_data_1[7]
port 19 nsew
flabel metal2 s 11610 14397 11666 15197 0 FreeSans 280 90 0 0 input_data_2[0]
port 20 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 input_data_2[1]
port 21 nsew
flabel metal3 s 12253 12248 13053 12368 0 FreeSans 600 0 0 0 input_data_2[2]
port 22 nsew
flabel metal2 s 2594 14397 2650 15197 0 FreeSans 280 90 0 0 input_data_2[3]
port 23 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 input_data_2[4]
port 24 nsew
flabel metal3 s 0 2728 800 2848 0 FreeSans 600 0 0 0 input_data_2[5]
port 25 nsew
flabel metal3 s 12253 8168 13053 8288 0 FreeSans 600 0 0 0 input_data_2[6]
port 26 nsew
flabel metal2 s 1306 14397 1362 15197 0 FreeSans 280 90 0 0 input_data_2[7]
port 27 nsew
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 input_data_3[0]
port 28 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 input_data_3[1]
port 29 nsew
flabel metal2 s 9034 14397 9090 15197 0 FreeSans 280 90 0 0 input_data_3[2]
port 30 nsew
flabel metal3 s 12253 4088 13053 4208 0 FreeSans 600 0 0 0 input_data_3[3]
port 31 nsew
flabel metal2 s 1306 0 1362 800 0 FreeSans 280 90 0 0 input_data_3[4]
port 32 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 input_data_3[5]
port 33 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 input_data_3[6]
port 34 nsew
flabel metal3 s 12253 5448 13053 5568 0 FreeSans 600 0 0 0 input_data_3[7]
port 35 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 output_data[0]
port 36 nsew
flabel metal3 s 12253 13608 13053 13728 0 FreeSans 600 0 0 0 output_data[1]
port 37 nsew
flabel metal2 s 12898 14397 12954 15197 0 FreeSans 280 90 0 0 output_data[2]
port 38 nsew
flabel metal2 s 3882 14397 3938 15197 0 FreeSans 280 90 0 0 output_data[3]
port 39 nsew
flabel metal2 s 5170 14397 5226 15197 0 FreeSans 280 90 0 0 output_data[4]
port 40 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 output_data[5]
port 41 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 output_data[6]
port 42 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 output_data[7]
port 43 nsew
flabel metal3 s 12253 6808 13053 6928 0 FreeSans 600 0 0 0 reset
port 44 nsew
<< properties >>
string FIXED_BBOX 0 0 13053 15197
<< end >>
