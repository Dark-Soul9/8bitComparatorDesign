VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Comparator
  CLASS BLOCK ;
  FOREIGN Comparator ;
  ORIGIN 0.000 0.000 ;
  SIZE 65.265 BY 75.985 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.280 58.600 59.580 60.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.680 59.580 47.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 32.760 59.580 34.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.840 59.580 21.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.110 10.640 56.710 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.655 10.640 43.255 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.200 10.640 29.800 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.745 10.640 16.345 62.800 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.280 55.300 59.580 56.900 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 42.380 59.580 43.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.460 59.580 31.060 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 16.540 59.580 18.140 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.810 10.640 53.410 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.355 10.640 39.955 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.900 10.640 26.500 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 11.445 10.640 13.045 62.800 ;
    END
  END VPWR
  PIN clk
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END clk
  PIN input_data_0[0]
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END input_data_0[0]
  PIN input_data_0[1]
    PORT
      LAYER met2 ;
        RECT 32.290 71.985 32.570 75.985 ;
    END
  END input_data_0[1]
  PIN input_data_0[2]
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END input_data_0[2]
  PIN input_data_0[3]
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END input_data_0[3]
  PIN input_data_0[4]
    PORT
      LAYER met3 ;
        RECT 61.265 6.840 65.265 7.440 ;
    END
  END input_data_0[4]
  PIN input_data_0[5]
    PORT
      LAYER met3 ;
        RECT 61.265 47.640 65.265 48.240 ;
    END
  END input_data_0[5]
  PIN input_data_0[6]
    PORT
      LAYER met2 ;
        RECT 0.090 71.985 0.370 75.985 ;
    END
  END input_data_0[6]
  PIN input_data_0[7]
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END input_data_0[7]
  PIN input_data_1[0]
    PORT
      LAYER met2 ;
        RECT 51.610 71.985 51.890 75.985 ;
    END
  END input_data_1[0]
  PIN input_data_1[1]
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END input_data_1[1]
  PIN input_data_1[2]
    PORT
      LAYER met3 ;
        RECT 61.265 54.440 65.265 55.040 ;
    END
  END input_data_1[2]
  PIN input_data_1[3]
    PORT
      LAYER met3 ;
        RECT 61.265 13.640 65.265 14.240 ;
    END
  END input_data_1[3]
  PIN input_data_1[4]
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END input_data_1[4]
  PIN input_data_1[5]
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END input_data_1[5]
  PIN input_data_1[6]
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END input_data_1[6]
  PIN input_data_1[7]
    PORT
      LAYER met2 ;
        RECT 38.730 71.985 39.010 75.985 ;
    END
  END input_data_1[7]
  PIN input_data_2[0]
    PORT
      LAYER met2 ;
        RECT 58.050 71.985 58.330 75.985 ;
    END
  END input_data_2[0]
  PIN input_data_2[1]
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END input_data_2[1]
  PIN input_data_2[2]
    PORT
      LAYER met3 ;
        RECT 61.265 61.240 65.265 61.840 ;
    END
  END input_data_2[2]
  PIN input_data_2[3]
    PORT
      LAYER met2 ;
        RECT 12.970 71.985 13.250 75.985 ;
    END
  END input_data_2[3]
  PIN input_data_2[4]
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END input_data_2[4]
  PIN input_data_2[5]
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END input_data_2[5]
  PIN input_data_2[6]
    PORT
      LAYER met3 ;
        RECT 61.265 40.840 65.265 41.440 ;
    END
  END input_data_2[6]
  PIN input_data_2[7]
    PORT
      LAYER met2 ;
        RECT 6.530 71.985 6.810 75.985 ;
    END
  END input_data_2[7]
  PIN input_data_3[0]
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END input_data_3[0]
  PIN input_data_3[1]
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END input_data_3[1]
  PIN input_data_3[2]
    PORT
      LAYER met2 ;
        RECT 45.170 71.985 45.450 75.985 ;
    END
  END input_data_3[2]
  PIN input_data_3[3]
    PORT
      LAYER met3 ;
        RECT 61.265 20.440 65.265 21.040 ;
    END
  END input_data_3[3]
  PIN input_data_3[4]
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END input_data_3[4]
  PIN input_data_3[5]
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END input_data_3[5]
  PIN input_data_3[6]
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END input_data_3[6]
  PIN input_data_3[7]
    PORT
      LAYER met3 ;
        RECT 61.265 27.240 65.265 27.840 ;
    END
  END input_data_3[7]
  PIN output_data[0]
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END output_data[0]
  PIN output_data[1]
    PORT
      LAYER met3 ;
        RECT 61.265 68.040 65.265 68.640 ;
    END
  END output_data[1]
  PIN output_data[2]
    PORT
      LAYER met2 ;
        RECT 64.490 71.985 64.770 75.985 ;
    END
  END output_data[2]
  PIN output_data[3]
    PORT
      LAYER met2 ;
        RECT 19.410 71.985 19.690 75.985 ;
    END
  END output_data[3]
  PIN output_data[4]
    PORT
      LAYER met2 ;
        RECT 25.850 71.985 26.130 75.985 ;
    END
  END output_data[4]
  PIN output_data[5]
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END output_data[5]
  PIN output_data[6]
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END output_data[6]
  PIN output_data[7]
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END output_data[7]
  PIN reset
    PORT
      LAYER met3 ;
        RECT 61.265 34.040 65.265 34.640 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 59.340 62.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 64.790 63.200 ;
      LAYER met2 ;
        RECT 0.650 71.705 6.250 72.490 ;
        RECT 7.090 71.705 12.690 72.490 ;
        RECT 13.530 71.705 19.130 72.490 ;
        RECT 19.970 71.705 25.570 72.490 ;
        RECT 26.410 71.705 32.010 72.490 ;
        RECT 32.850 71.705 38.450 72.490 ;
        RECT 39.290 71.705 44.890 72.490 ;
        RECT 45.730 71.705 51.330 72.490 ;
        RECT 52.170 71.705 57.770 72.490 ;
        RECT 58.610 71.705 64.210 72.490 ;
        RECT 0.100 4.280 64.760 71.705 ;
        RECT 0.650 4.000 6.250 4.280 ;
        RECT 7.090 4.000 12.690 4.280 ;
        RECT 13.530 4.000 19.130 4.280 ;
        RECT 19.970 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.010 4.280 ;
        RECT 32.850 4.000 38.450 4.280 ;
        RECT 39.290 4.000 44.890 4.280 ;
        RECT 45.730 4.000 51.330 4.280 ;
        RECT 52.170 4.000 57.770 4.280 ;
        RECT 58.610 4.000 64.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 67.640 60.865 68.505 ;
        RECT 4.000 62.240 61.265 67.640 ;
        RECT 4.400 60.840 60.865 62.240 ;
        RECT 4.000 55.440 61.265 60.840 ;
        RECT 4.400 54.040 60.865 55.440 ;
        RECT 4.000 48.640 61.265 54.040 ;
        RECT 4.400 47.240 60.865 48.640 ;
        RECT 4.000 41.840 61.265 47.240 ;
        RECT 4.400 40.440 60.865 41.840 ;
        RECT 4.000 35.040 61.265 40.440 ;
        RECT 4.400 33.640 60.865 35.040 ;
        RECT 4.000 28.240 61.265 33.640 ;
        RECT 4.400 26.840 60.865 28.240 ;
        RECT 4.000 21.440 61.265 26.840 ;
        RECT 4.400 20.040 60.865 21.440 ;
        RECT 4.000 14.640 61.265 20.040 ;
        RECT 4.400 13.240 60.865 14.640 ;
        RECT 4.000 7.840 61.265 13.240 ;
        RECT 4.400 6.975 60.865 7.840 ;
      LAYER met4 ;
        RECT 37.095 13.095 37.425 49.465 ;
  END
END Comparator
END LIBRARY

